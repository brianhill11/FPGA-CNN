`ifndef SOFTMAX_WITH_LOSS_TEST_H
`define SOFTMAX_WITH_LOSS_TEST_H
reg [31:0] test_input [40000];
reg [31:0] test_label [5000];
reg [31:0] test_output [5000];
initial begin
test_input[0:7] = '{32'hc2b396b3, 32'hc25023d4, 32'h4201d56e, 32'h41c7c297, 32'hc20fc999, 32'h4130133a, 32'hc2540616, 32'h42941b6f};
test_label[0] = '{32'hc25023d4};
test_output[0] = '{32'h42fc2d59};
/*############ DEBUG ############
test_input[0:7] = '{-89.794337838, -52.0349894359, 32.4584292302, 24.9700152718, -35.9468726419, 11.0046941298, -53.0059437905, 74.0535794014};
test_label[0] = '{-52.0349894359};
test_output[0] = '{126.088568837};
############ END DEBUG ############*/
test_input[8:15] = '{32'hc21b936f, 32'hc14826ee, 32'hc2a24141, 32'hc1de1817, 32'hc25c7cff, 32'h4292c216, 32'hc198b047, 32'hc2b64ae8};
test_label[1] = '{32'hc1de1817};
test_output[1] = '{32'h42ca481b};
/*############ DEBUG ############
test_input[8:15] = '{-38.8939784469, -12.5095039018, -81.1274470641, -27.7617620836, -55.1220677192, 73.3790706841, -19.0860733695, -91.1463004197};
test_label[1] = '{-27.7617620836};
test_output[1] = '{101.140832768};
############ END DEBUG ############*/
test_input[16:23] = '{32'hc1fc17dd, 32'h420d9f3c, 32'h42a2162a, 32'hc2a30145, 32'h422da8ab, 32'hc2ad087f, 32'h4282c34e, 32'h423f840b};
test_label[2] = '{32'hc2ad087f};
test_output[2] = '{32'h43278f55};
/*############ DEBUG ############
test_input[16:23] = '{-31.5116529328, 35.4055040754, 81.0432912975, -81.5024832633, 43.4147144174, -86.5165945903, 65.3814564659, 47.8789469151};
test_label[2] = '{-86.5165945903};
test_output[2] = '{167.559886046};
############ END DEBUG ############*/
test_input[24:31] = '{32'h4233df12, 32'hc298b589, 32'h4225884c, 32'hc28496fe, 32'hc28dbbf6, 32'hc2b12860, 32'h42ade654, 32'h42c4dcca};
test_label[3] = '{32'hc298b589};
test_output[3] = '{32'h432ec92a};
/*############ DEBUG ############
test_input[24:31] = '{44.9678418937, -76.354558961, 41.3831019686, -66.2949034573, -70.8671076641, -88.5788611872, 86.9498574502, 98.4312297522};
test_label[3] = '{-76.354558961};
test_output[3] = '{174.785799034};
############ END DEBUG ############*/
test_input[32:39] = '{32'h40d0ba1b, 32'h4234408a, 32'hc2bd6431, 32'h4195f821, 32'hc0d74f7a, 32'hc2515bad, 32'hc0bde248, 32'hc2ae55d9};
test_label[4] = '{32'hc0bde248};
test_output[4] = '{32'h424bfcd3};
/*############ DEBUG ############
test_input[32:39] = '{6.52271788842, 45.063025612, -94.6956881177, 18.7461560667, -6.72845154669, -52.3395266431, -5.9338722616, -87.1676691855};
test_label[4] = '{-5.9338722616};
test_output[4] = '{50.9968978736};
############ END DEBUG ############*/
test_input[40:47] = '{32'h423d0a71, 32'hc197fed7, 32'hc23bfec1, 32'hc183c7b3, 32'h4289cd0b, 32'hc2b58590, 32'h41a0b767, 32'h4188ede3};
test_label[5] = '{32'hc2b58590};
test_output[5] = '{32'h431fa94e};
/*############ DEBUG ############
test_input[40:47] = '{47.2601969947, -18.9994329118, -46.9987820931, -16.4725096596, 68.9004729773, -90.7608671655, 20.0895517604, 17.1161554362};
test_label[5] = '{-90.7608671655};
test_output[5] = '{159.661340143};
############ END DEBUG ############*/
test_input[48:55] = '{32'hc26fc9ca, 32'hc211c90a, 32'h4219ba59, 32'h425ddca5, 32'hc204085e, 32'h42782354, 32'hc28d6b87, 32'hc2ac280e};
test_label[6] = '{32'h425ddca5};
test_output[6] = '{32'h40d240f0};
/*############ DEBUG ############
test_input[48:55] = '{-59.9470612565, -36.4463274772, 38.4319795522, 55.4654735192, -33.0081700952, 62.0344982751, -70.7100137666, -86.0782281384};
test_label[6] = '{55.4654735192};
test_output[6] = '{6.57042693758};
############ END DEBUG ############*/
test_input[56:63] = '{32'hc20df4b0, 32'hc1892ce9, 32'hc0527636, 32'h412f7020, 32'hc0699383, 32'hc2541e10, 32'h4267d7ae, 32'hc2bc2a3e};
test_label[7] = '{32'h4267d7ae};
test_output[7] = '{32'h80000000};
/*############ DEBUG ############
test_input[56:63] = '{-35.4889538082, -17.146928353, -3.28846502654, 10.964873838, -3.64962843692, -53.0293581368, 57.9606231357, -94.0825041819};
test_label[7] = '{57.9606231357};
test_output[7] = '{-0.0};
############ END DEBUG ############*/
test_input[64:71] = '{32'h41d91ad0, 32'hc2b71c14, 32'hc2be8ea1, 32'hc2b5f1e1, 32'hc209979b, 32'hc2b1969f, 32'hc234ca21, 32'hc2b4bc85};
test_label[8] = '{32'h41d91ad0};
test_output[8] = '{32'h80000000};
/*############ DEBUG ############
test_input[64:71] = '{27.1380922832, -91.5548371963, -95.2785711421, -90.9724228601, -34.3980509595, -88.794183747, -45.1973928089, -90.3682015346};
test_label[8] = '{27.1380922832};
test_output[8] = '{-0.0};
############ END DEBUG ############*/
test_input[72:79] = '{32'h4287d739, 32'h42ae51b3, 32'hc1ac7e17, 32'h428da6a4, 32'h4283eba5, 32'hc29b5175, 32'hc2481002, 32'hc1b9f006};
test_label[9] = '{32'hc1ac7e17};
test_output[9] = '{32'h42d97138};
/*############ DEBUG ############
test_input[72:79] = '{67.9203582228, 87.1595654847, -21.5615680768, 70.8254708908, 65.9602454877, -77.6590992277, -50.0156314135, -23.2421983504};
test_label[9] = '{-21.5615680768};
test_output[9] = '{108.721133647};
############ END DEBUG ############*/
test_input[80:87] = '{32'hc281ad8c, 32'hc21491bd, 32'h422c839a, 32'hc18adf78, 32'hc21190a0, 32'h42248ea9, 32'h426f17d5, 32'hc22dfe0f};
test_label[10] = '{32'h426f17d5};
test_output[10] = '{32'h33902cba};
/*############ DEBUG ############
test_input[80:87] = '{-64.8389617049, -37.1423237018, 43.1285162705, -17.3591147623, -36.3912365915, 41.1393163595, 59.7732745009, -43.4981035087};
test_label[10] = '{59.7732745009};
test_output[10] = '{6.71365849913e-08};
############ END DEBUG ############*/
test_input[88:95] = '{32'h42c7018c, 32'hc2a96f75, 32'h4296fab8, 32'hc28d4320, 32'hc08649f7, 32'hc00775c3, 32'h42baf2a4, 32'h4238b82a};
test_label[11] = '{32'h42baf2a4};
test_output[11] = '{32'h40c10236};
/*############ DEBUG ############
test_input[88:95] = '{99.5030203922, -84.7176932578, 75.4896861255, -70.63110705, -4.19652891114, -2.11656254932, 93.4739050621, 46.1798493549};
test_label[11] = '{93.4739050621};
test_output[11] = '{6.0315200594};
############ END DEBUG ############*/
test_input[96:103] = '{32'h4104efc2, 32'hc2b4f101, 32'h41ff6cd3, 32'hc1e3519f, 32'hc2176a6c, 32'hc256aa8a, 32'h419ff791, 32'hc0e78bbd};
test_label[12] = '{32'hc1e3519f};
test_output[12] = '{32'h42715f3b};
/*############ DEBUG ############
test_input[96:103] = '{8.30853444899, -90.4707092919, 31.9281359367, -28.4148548868, -37.853927457, -53.6665406787, 19.9958815501, -7.2358080461};
test_label[12] = '{-28.4148548868};
test_output[12] = '{60.3429973984};
############ END DEBUG ############*/
test_input[104:111] = '{32'hc206ddb0, 32'h4260e8d9, 32'hc20372c5, 32'h4229be41, 32'hc2ab6484, 32'h41111627, 32'h42b36d9d, 32'hc1b23f20};
test_label[13] = '{32'h4229be41};
test_output[13] = '{32'h423d1cfa};
/*############ DEBUG ############
test_input[104:111] = '{-33.7164908099, 56.2273901665, -32.8620792848, 42.4357930008, -85.6963181986, 9.06790830446, 89.7140889361, -22.2808235458};
test_label[13] = '{42.4357930008};
test_output[13] = '{47.2782959352};
############ END DEBUG ############*/
test_input[112:119] = '{32'h41a0712a, 32'h420445d6, 32'hc2347dd9, 32'hc268755d, 32'h42be2644, 32'hc289d902, 32'h429e5641, 32'h42adb349};
test_label[14] = '{32'h429e5641};
test_output[14] = '{32'h417e812b};
/*############ DEBUG ############
test_input[112:119] = '{20.0552553227, 33.0681986168, -45.1228988589, -58.1146138422, 95.074735072, -68.923846057, 79.1684682004, 86.8501676285};
test_label[14] = '{79.1684682004};
test_output[14] = '{15.9065349475};
############ END DEBUG ############*/
test_input[120:127] = '{32'hc2b71ac9, 32'hc2828e00, 32'h41415c70, 32'h42089afc, 32'hc22a1f63, 32'h40f9c931, 32'h42794f27, 32'hc26527cc};
test_label[15] = '{32'h40f9c931};
test_output[15] = '{32'h425a1600};
/*############ DEBUG ############
test_input[120:127] = '{-91.5523138338, -65.2773433098, 12.0850675638, 34.151353429, -42.5306515863, 7.80580958683, 62.3272955061, -57.2888627938};
test_label[15] = '{7.80580958683};
test_output[15] = '{54.5214859193};
############ END DEBUG ############*/
test_input[128:135] = '{32'h42982f97, 32'hc27b9dbb, 32'h4298f5aa, 32'h4294f94a, 32'hc228e445, 32'h420a0187, 32'h42bb6516, 32'hc199b225};
test_label[16] = '{32'hc199b225};
test_output[16] = '{32'h42e1d1a0};
/*############ DEBUG ############
test_input[128:135] = '{76.092950564, -62.9040349921, 76.4798138911, 74.4868949147, -42.2229197668, 34.5014915675, 93.6974364935, -19.2119853486};
test_label[16] = '{-19.2119853486};
test_output[16] = '{112.909421902};
############ END DEBUG ############*/
test_input[136:143] = '{32'h416f0660, 32'h4213d1fd, 32'hc1a7c7ad, 32'h418b6d51, 32'h423ad850, 32'hc29278b5, 32'h422e0ed5, 32'hc1024d51};
test_label[17] = '{32'hc29278b5};
test_output[17] = '{32'h42eff96a};
/*############ DEBUG ############
test_input[136:143] = '{14.9390565042, 36.9550672354, -20.9724978261, 17.4283776701, 46.7112415114, -73.2357554403, 43.5144846112, -8.14387615104};
test_label[17] = '{-73.2357554403};
test_output[17] = '{119.987133159};
############ END DEBUG ############*/
test_input[144:151] = '{32'h418d4324, 32'h429c54bd, 32'h4221b6cd, 32'h42736e9d, 32'hc2beb0e1, 32'hc244fcf3, 32'hc2c1fbe7, 32'h42bc588d};
test_label[18] = '{32'hc2beb0e1};
test_output[18] = '{32'h433d84b7};
/*############ DEBUG ############
test_input[144:151] = '{17.6577827628, 78.1655067857, 40.4285145729, 60.8580203759, -95.3454654199, -49.2470200972, -96.9919960659, 94.1729525852};
test_label[18] = '{-95.3454654199};
test_output[18] = '{189.518418117};
############ END DEBUG ############*/
test_input[152:159] = '{32'hc25cf7c8, 32'hc1ffc2f4, 32'h41cd74ea, 32'hc29b58c1, 32'hc2b35333, 32'h428a8506, 32'hc2697874, 32'h404dfa50};
test_label[19] = '{32'hc2697874};
test_output[19] = '{32'h42ff4140};
/*############ DEBUG ############
test_input[152:159] = '{-55.2419734732, -31.9701928566, 25.682087357, -77.6733504992, -89.6624953566, 69.2598077937, -58.367629866, 3.21840296515};
test_label[19] = '{-58.367629866};
test_output[19] = '{127.62743766};
############ END DEBUG ############*/
test_input[160:167] = '{32'h41ee7ebd, 32'hc28e07c5, 32'hc29ddb57, 32'hc1eb5978, 32'h428d3aa0, 32'h4255f07d, 32'hc18021d7, 32'hc265865c};
test_label[20] = '{32'h41ee7ebd};
test_output[20] = '{32'h422335e3};
/*############ DEBUG ############
test_input[160:167] = '{29.811883093, -71.0151785609, -78.9283996049, -29.4186853031, 70.614505604, 53.4848514658, -16.0165229678, -57.3812095405};
test_label[20] = '{29.811883093};
test_output[20] = '{40.8026225474};
############ END DEBUG ############*/
test_input[168:175] = '{32'hc2b60383, 32'hc294e99a, 32'h41f8d3c7, 32'h4137a88d, 32'hc1253fd7, 32'hc2a10bbb, 32'hc2a4c289, 32'hc225f914};
test_label[21] = '{32'hc225f914};
test_output[21] = '{32'h4291317c};
/*############ DEBUG ############
test_input[168:175] = '{-91.0068565189, -74.4562499223, 31.1034070773, 11.4786500937, -10.3280855852, -80.5229092417, -82.3799533217, -41.4932415487};
test_label[21] = '{-41.4932415487};
test_output[21] = '{72.596648629};
############ END DEBUG ############*/
test_input[176:183] = '{32'hc0847bc2, 32'hc1295de0, 32'h42779bde, 32'h429f14b6, 32'hc2390b24, 32'hc166c80b, 32'hbf7b81eb, 32'h427d6f47};
test_label[22] = '{32'h429f14b6};
test_output[22] = '{32'h33f875c4};
/*############ DEBUG ############
test_input[176:183] = '{-4.14010692551, -10.5854184477, 61.9022122762, 79.5404500162, -46.2608791918, -14.4238383642, -0.982451117159, 63.358670279};
test_label[22] = '{79.5404500162};
test_output[22] = '{1.15698212154e-07};
############ END DEBUG ############*/
test_input[184:191] = '{32'hc274461f, 32'h4292b433, 32'hc2b9ddf2, 32'hc256df51, 32'h41810948, 32'hc1389924, 32'h428401fa, 32'h42685146};
test_label[23] = '{32'hc274461f};
test_output[23] = '{32'h43066bcc};
/*############ DEBUG ############
test_input[184:191] = '{-61.0684768049, 73.351953817, -92.9334899278, -53.7180819062, 16.1295311393, -11.5373877929, 66.0038606512, 58.0793704943};
test_label[23] = '{-61.0684768049};
test_output[23] = '{134.421074466};
############ END DEBUG ############*/
test_input[192:199] = '{32'h41d64bb8, 32'hc28ab58f, 32'h41c4a044, 32'hc2518c64, 32'h4169c769, 32'hc2ab9436, 32'hc22bc8b9, 32'hc2bb8a26};
test_label[24] = '{32'hc22bc8b9};
test_output[24] = '{32'h428baca7};
/*############ DEBUG ############
test_input[192:199] = '{26.7869718162, -69.35460866, 24.5782541381, -52.3870990162, 14.6111843809, -85.789472338, -42.9460186341, -93.7698234025};
test_label[24] = '{-42.9460186341};
test_output[24] = '{69.8372122255};
############ END DEBUG ############*/
test_input[200:207] = '{32'hc239b6f7, 32'h420aeb29, 32'h4162b290, 32'h403a3a53, 32'hc03a68dc, 32'h42bbb303, 32'hc1bf479a, 32'hc0aad3f8};
test_label[25] = '{32'hc03a68dc};
test_output[25] = '{32'h42c1864a};
/*############ DEBUG ############
test_input[200:207] = '{-46.4286776974, 34.7296504282, 14.1685947571, 2.90980980641, -2.91265006897, 93.8496340176, -23.9099618475, -5.33837498709};
test_label[25] = '{-2.91265006897};
test_output[25] = '{96.7622840865};
############ END DEBUG ############*/
test_input[208:215] = '{32'hc26232d7, 32'hc2ab58b1, 32'hc2804470, 32'hc19057bd, 32'hc234bb34, 32'hc283a66a, 32'hc1fd8b43, 32'h4281c6d0};
test_label[26] = '{32'hc2804470};
test_output[26] = '{32'h430105a0};
/*############ DEBUG ############
test_input[208:215] = '{-56.549647373, -85.6732269431, -64.1336650649, -18.0428417514, -45.1828166849, -65.8250271204, -31.6929986514, 64.8883053218};
test_label[26] = '{-64.1336650649};
test_output[26] = '{129.021970387};
############ END DEBUG ############*/
test_input[216:223] = '{32'h41f15a07, 32'h42955801, 32'h41c59d4f, 32'h42b705f5, 32'h426bfa39, 32'hc2c05c70, 32'h429b5577, 32'hc2ae02f4};
test_label[27] = '{32'h42b705f5};
test_output[27] = '{32'h3588e0af};
/*############ DEBUG ############
test_input[216:223] = '{30.1689589797, 74.6718825365, 24.7018115563, 91.5116324615, 58.9943587567, -96.1805400137, 77.666923588, -87.0057663392};
test_label[27] = '{91.5116324615};
test_output[27] = '{1.01981809407e-06};
############ END DEBUG ############*/
test_input[224:231] = '{32'hc23a90c2, 32'hc27b05c3, 32'hc2af42dd, 32'h4008625f, 32'h42aec16e, 32'hc112974d, 32'hc29ef9bc, 32'hc23174dd};
test_label[28] = '{32'h4008625f};
test_output[28] = '{32'h42aa7e5b};
/*############ DEBUG ############
test_input[224:231] = '{-46.6413656239, -62.7556284365, -87.6305888044, 2.13100414137, 87.3777901931, -9.16193872166, -79.4877630402, -44.364124369};
test_label[28] = '{2.13100414137};
test_output[28] = '{85.2467860517};
############ END DEBUG ############*/
test_input[232:239] = '{32'hc21455ba, 32'h40c63449, 32'h42b0f554, 32'h40ba50f7, 32'hc18aea72, 32'h419e84bd, 32'h42b9a751, 32'h41b5fedb};
test_label[29] = '{32'h40ba50f7};
test_output[29] = '{32'h42ae08d6};
/*############ DEBUG ############
test_input[232:239] = '{-37.0837156105, 6.19388228594, 88.4791538801, 5.82238323007, -17.3644753364, 19.8148145068, 92.8267868219, 22.7494409561};
test_label[29] = '{5.82238323007};
test_output[29] = '{87.0172580185};
############ END DEBUG ############*/
test_input[240:247] = '{32'h42943b44, 32'hc2baad43, 32'hc1d75663, 32'h42a4b59e, 32'h41be1c4a, 32'hc1e540f9, 32'h40de1554, 32'h423dbe3d};
test_label[30] = '{32'hc1e540f9};
test_output[30] = '{32'h42de05ff};
/*############ DEBUG ############
test_input[240:247] = '{74.1157513746, -93.3384034778, -26.9171808739, 82.3547238115, 23.7638135063, -28.6567241066, 6.94010350457, 47.4357804042};
test_label[30] = '{-28.6567241066};
test_output[30] = '{111.011712039};
############ END DEBUG ############*/
test_input[248:255] = '{32'hc266df26, 32'h42bcfcb5, 32'hc154911d, 32'h42a73799, 32'hc1f57ec2, 32'h41d05ea4, 32'hc2605af5, 32'h41a3b998};
test_label[31] = '{32'h42a73799};
test_output[31] = '{32'h412e28f8};
/*############ DEBUG ############
test_input[248:255] = '{-57.7179177092, 94.4935707846, -13.2854284037, 83.6085869191, -30.6868935498, 26.046210942, -56.0888262048, 20.465621829};
test_label[31] = '{83.6085869191};
test_output[31] = '{10.8850026028};
############ END DEBUG ############*/
test_input[256:263] = '{32'hc1336ea8, 32'hc0e9b269, 32'h42968da1, 32'h42458643, 32'h420845ef, 32'hc13ac14d, 32'h41e8caf3, 32'h412b7f3a};
test_label[32] = '{32'hc0e9b269};
test_output[32] = '{32'h42a528c8};
/*############ DEBUG ############
test_input[256:263] = '{-11.2145154906, -7.30302881084, 75.2766201236, 49.3811157441, 34.0682926198, -11.6721922274, 29.0990964767, 10.7185612418};
test_label[32] = '{-7.30302881084};
test_output[32] = '{82.5796489345};
############ END DEBUG ############*/
test_input[264:271] = '{32'h421b64a9, 32'hc2c3d566, 32'h424b2215, 32'h42399060, 32'h42911cce, 32'hc206520b, 32'hc26130ad, 32'hc2528c6f};
test_label[33] = '{32'hc206520b};
test_output[33] = '{32'h42d445d4};
/*############ DEBUG ############
test_input[264:271] = '{38.8483017843, -97.9167901174, 50.783283767, 46.3909904902, 72.5562620674, -33.5801197595, -56.2975361514, -52.6371426773};
test_label[33] = '{-33.5801197595};
test_output[33] = '{106.136381827};
############ END DEBUG ############*/
test_input[272:279] = '{32'hc28e9a8c, 32'hc299eb5e, 32'hc0e3b89f, 32'hc2c1552e, 32'h42801fea, 32'hc23b5951, 32'hc006fd1c, 32'h421ec981};
test_label[34] = '{32'hc2c1552e};
test_output[34] = '{32'h4320ba8c};
/*############ DEBUG ############
test_input[272:279] = '{-71.3018467472, -76.959704765, -7.11628676602, -96.6663689555, 64.0623324841, -46.8372221405, -2.10919849941, 39.6967807411};
test_label[34] = '{-96.6663689555};
test_output[34] = '{160.72870144};
############ END DEBUG ############*/
test_input[280:287] = '{32'hc20a90a4, 32'hc20a5e06, 32'h41e9a8dd, 32'hc0c53373, 32'hc1db600c, 32'h4102df31, 32'hc2460947, 32'hc28a8804};
test_label[35] = '{32'hc28a8804};
test_output[35] = '{32'h42c4f23c};
/*############ DEBUG ############
test_input[280:287] = '{-34.6412501712, -34.5918199352, 29.207453178, -6.16253036598, -27.4218976475, 8.17948978419, -49.5090602557, -69.2656591829};
test_label[35] = '{-69.2656591829};
test_output[35] = '{98.4731123617};
############ END DEBUG ############*/
test_input[288:295] = '{32'hc288f5fa, 32'h428f81a7, 32'h42b418d3, 32'h3ec371c2, 32'hc20215f7, 32'hc26a3a96, 32'h42c06c6f, 32'h4175d88b};
test_label[36] = '{32'hc20215f7};
test_output[36] = '{32'h4300bc3f};
/*############ DEBUG ############
test_input[288:295] = '{-68.4804214547, 71.753229472, 90.0484864102, 0.381727281471, -32.5214499524, -58.5572140225, 96.2117880866, 15.3653664923};
test_label[36] = '{-32.5214499524};
test_output[36] = '{128.735341117};
############ END DEBUG ############*/
test_input[296:303] = '{32'hc2889975, 32'h42c0742e, 32'h416a8529, 32'h42bdeb0e, 32'hc2af3901, 32'h42bb78a8, 32'hc1317053, 32'h427f9fd8};
test_label[37] = '{32'h416a8529};
test_output[37] = '{32'h42a3c290};
/*############ DEBUG ############
test_input[296:303] = '{-68.2997195456, 96.2269108856, 14.6575093413, 94.9590942454, -87.6113362397, 93.7356596051, -11.0899231065, 63.9060972977};
test_label[37] = '{14.6575093413};
test_output[37] = '{81.8800076438};
############ END DEBUG ############*/
test_input[304:311] = '{32'hc1beab51, 32'hc2576e82, 32'hc1b6ae5c, 32'hc286f74e, 32'h42acfa47, 32'hc2151c86, 32'h41f0d929, 32'h42868c86};
test_label[38] = '{32'hc1b6ae5c};
test_output[38] = '{32'h42daa5de};
/*############ DEBUG ############
test_input[304:311] = '{-23.8336513097, -53.8579186141, -22.8351369198, -67.4830190574, 86.4888215334, -37.2778544381, 30.1060356114, 67.2744632474};
test_label[38] = '{-22.8351369198};
test_output[38] = '{109.323958458};
############ END DEBUG ############*/
test_input[312:319] = '{32'hc29cfb04, 32'hc1a818ce, 32'h42853f95, 32'h42bc9004, 32'hc235a473, 32'h4241c166, 32'h40881611, 32'hc1775d61};
test_label[39] = '{32'hc1775d61};
test_output[39] = '{32'h42db7bb0};
/*############ DEBUG ############
test_input[312:319] = '{-78.4902657858, -21.0121113346, 66.6241836494, 94.2812770031, -45.4105934017, 48.4388661315, 4.25269355245, -15.4602978287};
test_label[39] = '{-15.4602978287};
test_output[39] = '{109.741574832};
############ END DEBUG ############*/
test_input[320:327] = '{32'h421c4793, 32'h42a1cd55, 32'h420a1f65, 32'h42809ac6, 32'hc2bb0188, 32'hc22fde3e, 32'hc28d470f, 32'hc2829d18};
test_label[40] = '{32'h420a1f65};
test_output[40] = '{32'h42397b46};
/*############ DEBUG ############
test_input[320:327] = '{39.0698968603, 80.9010404656, 34.5306575723, 64.3022882938, -93.5029890671, -43.9670332474, -70.6387845728, -65.3068208851};
test_label[40] = '{34.5306575723};
test_output[40] = '{46.3703829551};
############ END DEBUG ############*/
test_input[328:335] = '{32'hc1d04d75, 32'h42abe13b, 32'h401e6822, 32'h4240e398, 32'h41fababa, 32'h417d5559, 32'hc20e65da, 32'h42b4dca9};
test_label[41] = '{32'h41fababa};
test_output[41] = '{32'h426c675f};
/*############ DEBUG ############
test_input[328:335] = '{-26.0378206866, 85.9399012009, 2.4751057718, 48.2222591297, 31.3411753125, 15.833336611, -35.5994656189, 90.4309762541};
test_label[41] = '{31.3411753125};
test_output[41] = '{59.1009471783};
############ END DEBUG ############*/
test_input[336:343] = '{32'hc28512df, 32'h4214b7ac, 32'h428e1eda, 32'hc27144b5, 32'h42952b21, 32'hc2baa0cc, 32'h41694010, 32'hc23411bb};
test_label[42] = '{32'hc28512df};
test_output[42] = '{32'h430d2670};
/*############ DEBUG ############
test_input[336:343] = '{-66.536854816, 37.1793677561, 71.0602532841, -60.3170952607, 74.5842348381, -93.3140555496, 14.578140425, -45.0173152703};
test_label[42] = '{-66.536854816};
test_output[42] = '{141.15014524};
############ END DEBUG ############*/
test_input[344:351] = '{32'h41a8272d, 32'hc23fcd39, 32'hc29627be, 32'h40ab6f09, 32'h428ce82b, 32'hc29d4f06, 32'hc29b959b, 32'h42ac0eaa};
test_label[43] = '{32'h40ab6f09};
test_output[43] = '{32'h42a157b9};
/*############ DEBUG ############
test_input[344:351] = '{21.0191278973, -47.9504136892, -75.0776240219, 5.35730421401, 70.4534562548, -78.6543429671, -77.7921955634, 86.0286391118};
test_label[43] = '{5.35730421401};
test_output[43] = '{80.6713350699};
############ END DEBUG ############*/
test_input[352:359] = '{32'hc20c660d, 32'h422ef5c4, 32'hc2ad3f14, 32'h42929842, 32'hc2b4a400, 32'h42adce60, 32'h418ca5d7, 32'hc28e7bdc};
test_label[44] = '{32'hc28e7bdc};
test_output[44] = '{32'h431e251e};
/*############ DEBUG ############
test_input[352:359] = '{-35.0996607867, 43.7400067595, -86.6231959365, 73.2973780075, -90.3203137033, 86.9030789963, 17.5809756037, -71.2419117293};
test_label[44] = '{-71.2419117293};
test_output[44] = '{158.144991959};
############ END DEBUG ############*/
test_input[360:367] = '{32'hc283fc9d, 32'h427c5049, 32'h42ab73e1, 32'hc175d92d, 32'h4264e1e9, 32'hc29b6d0c, 32'h42357a50, 32'hc1dc8f1c};
test_label[45] = '{32'hc1dc8f1c};
test_output[45] = '{32'h42e297a8};
/*############ DEBUG ############
test_input[360:367] = '{-65.9933829554, 63.078402756, 85.7263279475, -15.3655217351, 57.2206146533, -77.7129783935, 45.3694457368, -27.5698774439};
test_label[45] = '{-27.5698774439};
test_output[45] = '{113.296205392};
############ END DEBUG ############*/
test_input[368:375] = '{32'h4222b8d7, 32'hc1e66125, 32'h41e9ae63, 32'hc141f00b, 32'hc28fed6c, 32'h428c3b63, 32'h420e8508, 32'hc282caed};
test_label[46] = '{32'hc1e66125};
test_output[46] = '{32'h42c5d3ac};
/*############ DEBUG ############
test_input[368:375] = '{40.6805079489, -28.7974346312, 29.2101495056, -12.1211042958, -71.9637154125, 70.1159862908, 35.6299150984, -65.3963405996};
test_label[46] = '{-28.7974346312};
test_output[46] = '{98.913420922};
############ END DEBUG ############*/
test_input[376:383] = '{32'hc1be6142, 32'hc1976d74, 32'h4276568b, 32'hc1df8be6, 32'hc25b4ac4, 32'h40e1e339, 32'hc1ecc27e, 32'hc211911d};
test_label[47] = '{32'hc1be6142};
test_output[47] = '{32'h42aac396};
/*############ DEBUG ############
test_input[376:383] = '{-23.7974889657, -18.9284437891, 61.5845135945, -27.9433103336, -54.8230141742, 7.0589869215, -29.5949672414, -36.3917113209};
test_label[47] = '{-23.7974889657};
test_output[47] = '{85.3820025602};
############ END DEBUG ############*/
test_input[384:391] = '{32'hc1ad9a16, 32'h428f6c61, 32'h425257fb, 32'hc2690afa, 32'hc2be00d9, 32'hc2a2f25d, 32'h425335f0, 32'h406905b1};
test_label[48] = '{32'h428f6c61};
test_output[48] = '{32'h323e4e3a};
/*############ DEBUG ############
test_input[384:391] = '{-21.7002364793, 71.7116779821, 52.585920202, -58.2607188185, -95.0016587533, -81.4733660463, 52.8026727636, 3.64097242296};
test_label[48] = '{71.7116779821};
test_output[48] = '{1.10772421849e-08};
############ END DEBUG ############*/
test_input[392:399] = '{32'h3f358714, 32'hc257c004, 32'hc19dcfec, 32'h42b358f8, 32'h408b45e9, 32'h4254017a, 32'hc0667377, 32'hc258bd2d};
test_label[49] = '{32'hc257c004};
test_output[49] = '{32'h430f9c7d};
/*############ DEBUG ############
test_input[392:399] = '{0.709092357467, -53.9375169953, -19.7265235152, 89.6737690632, 4.35228418823, 53.0014426353, -3.60079740671, -54.1847426903};
test_label[49] = '{-53.9375169953};
test_output[49] = '{143.611286058};
############ END DEBUG ############*/
test_input[400:407] = '{32'hc2b8247d, 32'hc2b87909, 32'h40d25c51, 32'hbc78d063, 32'h41b4f248, 32'hc23f6651, 32'h42bb9ca1, 32'hc1c12abe};
test_label[50] = '{32'h41b4f248};
test_output[50] = '{32'h428e600f};
/*############ DEBUG ############
test_input[400:407] = '{-92.0712691509, -92.2363988946, 6.57376897447, -0.0151864017586, 22.6183006812, -47.8499168855, 93.8059144661, -24.1458710589};
test_label[50] = '{22.6183006812};
test_output[50] = '{71.187613785};
############ END DEBUG ############*/
test_input[408:415] = '{32'hc25a7216, 32'h422da5c6, 32'h42417c58, 32'hc13bceb8, 32'h406a5b95, 32'h40496fbc, 32'hc2923dab, 32'h42b88c5b};
test_label[51] = '{32'h42417c58};
test_output[51] = '{32'h422f9c5e};
/*############ DEBUG ############
test_input[408:415] = '{-54.6114110172, 43.4118864629, 48.3714294827, -11.7379680504, 3.66183963716, 3.14744471775, -73.1204482728, 92.2741329751};
test_label[51] = '{48.3714294827};
test_output[51] = '{43.9027034925};
############ END DEBUG ############*/
test_input[416:423] = '{32'h42184f5e, 32'h429cfd11, 32'h4282ec08, 32'hc2b449b0, 32'hc2b0327b, 32'h4110266c, 32'h42a565d7, 32'h414a1491};
test_label[52] = '{32'h4282ec08};
test_output[52] = '{32'h418a0593};
/*############ DEBUG ############
test_input[416:423] = '{38.0775054054, 78.4942738784, 65.461002024, -90.1439245384, -88.0985957443, 9.00937995514, 82.6989085678, 12.6300209871};
test_label[52] = '{65.461002024};
test_output[52] = '{17.2527225137};
############ END DEBUG ############*/
test_input[424:431] = '{32'h4299f7cf, 32'h42ab26a1, 32'hc25265d4, 32'hc2019546, 32'h4236f2cb, 32'hc02bda04, 32'h41c9eced, 32'h40db3ef0};
test_label[53] = '{32'h41c9eced};
test_output[53] = '{32'h427156fc};
/*############ DEBUG ############
test_input[424:431] = '{76.9840033319, 85.5754452816, -52.5994417529, -32.3957752635, 45.7371019914, -2.68518151218, 25.240685884, 6.85143280327};
test_label[53] = '{25.240685884};
test_output[53] = '{60.3349450685};
############ END DEBUG ############*/
test_input[432:439] = '{32'h42bd5f85, 32'h41068304, 32'hc2c0193a, 32'hc2812160, 32'hc2957020, 32'h4175215c, 32'hc09ff843, 32'h41283fed};
test_label[54] = '{32'h41068304};
test_output[54] = '{32'h42ac8f24};
/*############ DEBUG ############
test_input[432:439] = '{94.6865600211, 8.406986371, -96.0492739484, -64.565184224, -74.7189956341, 15.3206440357, -4.99905537354, 10.5156067226};
test_label[54] = '{8.406986371};
test_output[54] = '{86.2795736501};
############ END DEBUG ############*/
test_input[440:447] = '{32'hc22fa1ed, 32'h4166be32, 32'hc13c2154, 32'hc28bb852, 32'hc1c00aca, 32'hc2a9f4f3, 32'h429fc99d, 32'h421ab72a};
test_label[55] = '{32'h429fc99d};
test_output[55] = '{32'h80000000};
/*############ DEBUG ############
test_input[440:447] = '{-43.9081312207, 14.4214341213, -11.7581369227, -69.8599969661, -24.0052677767, -84.9784161873, 79.8937790307, 38.6788699627};
test_label[55] = '{79.8937790307};
test_output[55] = '{-0.0};
############ END DEBUG ############*/
test_input[448:455] = '{32'h42630970, 32'h42245306, 32'hc25dc909, 32'hc13127b3, 32'hc2b9b18a, 32'hc24e5de4, 32'h41f0ba97, 32'hc156424a};
test_label[56] = '{32'hc2b9b18a};
test_output[56] = '{32'h43159b21};
/*############ DEBUG ############
test_input[448:455] = '{56.7592147614, 41.0810793413, -55.4463246234, -11.0721918048, -92.846758545, -51.5916919655, 30.0911092296, -13.391184244};
test_label[56] = '{-92.846758545};
test_output[56] = '{149.605973462};
############ END DEBUG ############*/
test_input[456:463] = '{32'h4289f12f, 32'hc250dcbe, 32'h3ffac3ad, 32'hc220edc5, 32'hc1a9cbfb, 32'h42a84bcd, 32'h4205b517, 32'h42bb8a98};
test_label[57] = '{32'hc220edc5};
test_output[57] = '{32'h430600c1};
/*############ DEBUG ############
test_input[456:463] = '{68.971065032, -52.2155669036, 1.95909653766, -40.2321961394, -21.224599667, 84.1480504356, 33.4268472907, 93.7706880834};
test_label[57] = '{-40.2321961394};
test_output[57] = '{134.002950433};
############ END DEBUG ############*/
test_input[464:471] = '{32'h418d7c6d, 32'hc1bddb73, 32'h422881a5, 32'h42b46726, 32'h4034d518, 32'hc2a1b30f, 32'hc23a69e9, 32'hc1c7df5c};
test_label[58] = '{32'hc2a1b30f};
test_output[58] = '{32'h432b0d1a};
/*############ DEBUG ############
test_input[464:471] = '{17.6857544991, -23.7321533827, 42.1266051227, 90.2014631738, 2.82550611427, -80.8497208878, -46.6034283148, -24.9840630322};
test_label[58] = '{-80.8497208878};
test_output[58] = '{171.051184062};
############ END DEBUG ############*/
test_input[472:479] = '{32'h42522195, 32'h4259c933, 32'h42c08b5e, 32'hc23ddf92, 32'hc2ad3805, 32'hc2794ebf, 32'h42c159e8, 32'h4266a575};
test_label[59] = '{32'h4266a575};
test_output[59] = '{32'h421e1a4a};
/*############ DEBUG ############
test_input[472:479] = '{52.5327946737, 54.44648412, 96.2722036109, -47.4683307626, -86.6094132323, -62.3269016256, 96.675599178, 57.6615808047};
test_label[59] = '{57.6615808047};
test_output[59] = '{39.5256723275};
############ END DEBUG ############*/
test_input[480:487] = '{32'h425cbc83, 32'h4170a4b1, 32'h420c742b, 32'hc1addb35, 32'hc23a2828, 32'hc1a01179, 32'hc28b0b01, 32'h4238a1a6};
test_label[60] = '{32'hc1addb35};
test_output[60] = '{32'h4299d51f};
/*############ DEBUG ############
test_input[480:487] = '{55.1840946989, 15.0402078833, 35.1134468019, -21.7320340649, -46.5392145046, -20.0085317695, -69.5214944211, 46.1578582592};
test_label[60] = '{-21.7320340649};
test_output[60] = '{76.9162489725};
############ END DEBUG ############*/
test_input[488:495] = '{32'h41f34f21, 32'h422cdc13, 32'h425ef539, 32'h42211628, 32'hc20f3abb, 32'h40536e1b, 32'h40ed4f50, 32'h42437cda};
test_label[61] = '{32'h41f34f21};
test_output[61] = '{32'h41ca9d75};
/*############ DEBUG ############
test_input[488:495] = '{30.4136362382, 43.214914568, 55.7394758412, 40.2716375504, -35.80735252, 3.30359530021, 7.41593177903, 48.8719243332};
test_label[61] = '{30.4136362382};
test_output[61] = '{25.3268839082};
############ END DEBUG ############*/
test_input[496:503] = '{32'h4222ff64, 32'hc1424041, 32'h425f9474, 32'h407d118c, 32'hc28943e1, 32'h42c5409f, 32'h42bc7928, 32'hc24ae0d0};
test_label[62] = '{32'hc28943e1};
test_output[62] = '{32'h43274568};
/*############ DEBUG ############
test_input[496:503] = '{40.7494031861, -12.1406865269, 55.8949718499, 3.95419592788, -68.6325761247, 98.626216652, 94.2366330807, -50.7195452243};
test_label[62] = '{-68.6325761247};
test_output[62] = '{167.271122348};
############ END DEBUG ############*/
test_input[504:511] = '{32'hc2b66d4a, 32'hc29175f0, 32'hc2c6c84f, 32'h42b343da, 32'h42c6891c, 32'h412dc3ad, 32'hc1ba9137, 32'hc235cfb6};
test_label[63] = '{32'h42b343da};
test_output[63] = '{32'h411a2a53};
/*############ DEBUG ############
test_input[504:511] = '{-91.2134545739, -72.7303460415, -99.3912266847, 89.6325224517, 99.2677898072, 10.8602727016, -23.3209063778, -45.4528440413};
test_label[63] = '{89.6325224517};
test_output[63] = '{9.63533273511};
############ END DEBUG ############*/
test_input[512:519] = '{32'hc24ebfd6, 32'h429758ad, 32'h422f0a1d, 32'hc2a70955, 32'h42b2d2da, 32'h426e8813, 32'hbf33db67, 32'hc2c655cd};
test_label[64] = '{32'h429758ad};
test_output[64] = '{32'h415bd168};
/*############ DEBUG ############
test_input[512:519] = '{-51.6873400294, 75.6731966399, 43.7598764504, -83.5182244186, 89.4118206041, 59.6328863039, -0.70256655085, -99.1675779809};
test_label[64] = '{75.6731966399};
test_output[64] = '{13.7386250441};
############ END DEBUG ############*/
test_input[520:527] = '{32'h41f05d07, 32'h421f7374, 32'h42991f05, 32'h4257999a, 32'h428ccf93, 32'h42032c44, 32'h422ecbbe, 32'h4298c6e3};
test_label[65] = '{32'h421f7374};
test_output[65] = '{32'h42153d34};
/*############ DEBUG ############
test_input[520:527] = '{30.0454240488, 39.8627453218, 76.5605831761, 53.9000019444, 70.405421058, 32.7932269415, 43.6989688119, 76.3884493682};
test_label[65] = '{39.8627453218};
test_output[65] = '{37.3097690219};
############ END DEBUG ############*/
test_input[528:535] = '{32'h42aeafd1, 32'h424c56fb, 32'h42c56b60, 32'hc25dcf84, 32'hc202910c, 32'hc1fbedef, 32'hc19d3cd5, 32'h41bc7b15};
test_label[66] = '{32'hc202910c};
test_output[66] = '{32'h430359f4};
/*############ DEBUG ############
test_input[528:535] = '{87.3433941076, 51.0849432977, 98.7097189464, -55.452652517, -32.6416478536, -31.4911784183, -19.6547023417, 23.5600990891};
test_label[66] = '{-32.6416478536};
test_output[66] = '{131.351378379};
############ END DEBUG ############*/
test_input[536:543] = '{32'hc16e6376, 32'hc2660010, 32'hbf3ab7aa, 32'hc2abb8e6, 32'h41f79ad9, 32'h42acc681, 32'hc2bc822b, 32'h4278e824};
test_label[67] = '{32'hc2bc822b};
test_output[67] = '{32'h4334a456};
/*############ DEBUG ############
test_input[536:543] = '{-14.8992820955, -57.500060958, -0.729364996124, -85.8611307736, 30.9506086172, 86.3877033243, -94.2542305493, 62.2266994937};
test_label[67] = '{-94.2542305493};
test_output[67] = '{180.641933874};
############ END DEBUG ############*/
test_input[544:551] = '{32'hc147fec5, 32'h426be22d, 32'h4271d168, 32'h426d7469, 32'h41798b3b, 32'h41d3cbb3, 32'hc2300f93, 32'hc25e28ec};
test_label[68] = '{32'h4271d168};
test_output[68] = '{32'h3ee49550};
/*############ DEBUG ############
test_input[544:551] = '{-12.4996996027, 58.9708746373, 60.4544977284, 59.3636830556, 15.5964915929, 26.474462334, -44.0152097597, -55.5399618207};
test_label[68] = '{60.4544977284};
test_output[68] = '{0.446451650618};
############ END DEBUG ############*/
test_input[552:559] = '{32'h41b0d11d, 32'h417d2a0a, 32'hc2818dc4, 32'h4285da4c, 32'hc09a047d, 32'h42b2f73f, 32'h42070261, 32'h42a27d4e};
test_label[69] = '{32'h4285da4c};
test_output[69] = '{32'h41b47457};
/*############ DEBUG ############
test_input[552:559] = '{22.1021062373, 15.8227630413, -64.7768870174, 66.9263623563, -4.81304773159, 89.4829040761, 33.7523237669, 81.2447386372};
test_label[69] = '{66.9263623563};
test_output[69] = '{22.5568060539};
############ END DEBUG ############*/
test_input[560:567] = '{32'h42866a05, 32'h42c418d1, 32'h417c0c95, 32'hc2be75f7, 32'hc1e84f0e, 32'hc1bed3f2, 32'h422bb865, 32'h4240617f};
test_label[70] = '{32'h42866a05};
test_output[70] = '{32'h41f6bb2f};
/*############ DEBUG ############
test_input[560:567] = '{67.2070689103, 98.0484668021, 15.7530715464, -95.2304003452, -29.0386012148, -23.8534893588, 42.930073567, 48.0952113787};
test_label[70] = '{67.2070689103};
test_output[70] = '{30.8413978918};
############ END DEBUG ############*/
test_input[568:575] = '{32'hc24974e7, 32'h41e00060, 32'h42bb76f4, 32'h4269c6af, 32'hc101181e, 32'hc18e094f, 32'hc21d3ea0, 32'h412eeca5};
test_label[71] = '{32'hc21d3ea0};
test_output[71] = '{32'h43050b22};
/*############ DEBUG ############
test_input[568:575] = '{-50.3641624162, 28.0001825618, 93.7323283558, 58.4440283293, -8.06838803344, -17.7545460541, -39.3111561616, 10.9327740808};
test_label[71] = '{-39.3111561616};
test_output[71] = '{133.043484517};
############ END DEBUG ############*/
test_input[576:583] = '{32'hc28efd7b, 32'hc234fc5a, 32'hc2816c87, 32'hc2883f5a, 32'h42a34738, 32'hc247e528, 32'h40b0f5ee, 32'h42a93b98};
test_label[72] = '{32'h40b0f5ee};
test_output[72] = '{32'h429e45a8};
/*############ DEBUG ############
test_input[576:583] = '{-71.4950785317, -45.2464377361, -64.7119637299, -68.1237329328, 81.6390981772, -49.9737845358, 5.53002063185, 84.6163943673};
test_label[72] = '{5.53002063185};
test_output[72] = '{79.1360495586};
############ END DEBUG ############*/
test_input[584:591] = '{32'hc26d5902, 32'h41e3f830, 32'hc1c1edcb, 32'h41bf593b, 32'h429a6dfd, 32'h428e7829, 32'h42a46331, 32'h42868433};
test_label[73] = '{32'h42868433};
test_output[73] = '{32'h416f141c};
/*############ DEBUG ############
test_input[584:591] = '{-59.3369217324, 28.4961846462, -24.2411095971, 23.9185686592, 77.2148214506, 71.2346913144, 82.1937360228, 67.2582021473};
test_label[73] = '{67.2582021473};
test_output[73] = '{14.9424094387};
############ END DEBUG ############*/
test_input[592:599] = '{32'hc20a33bf, 32'hc24fb541, 32'h42c69b9d, 32'hc2bcb1c9, 32'hc23ab9ef, 32'hc2ae9f85, 32'h402e5314, 32'h42178c5e};
test_label[74] = '{32'h402e5314};
test_output[74] = '{32'h42c12904};
/*############ DEBUG ############
test_input[592:599] = '{-34.5505346633, -51.9270072777, 99.3039312915, -94.3472372677, -46.6815768624, -87.3115615983, 2.72382071352, 37.8870764121};
test_label[74] = '{2.72382071352};
test_output[74] = '{96.580110578};
############ END DEBUG ############*/
test_input[600:607] = '{32'hc2873e1c, 32'h41578ee2, 32'h4218ad0f, 32'h4242ce4e, 32'h41b5ad79, 32'hc2248faa, 32'hc1ac74e0, 32'hc2303390};
test_label[75] = '{32'h4242ce4e};
test_output[75] = '{32'h37df9c4b};
/*############ DEBUG ############
test_input[600:607] = '{-67.6213099803, 13.4723839529, 38.169002705, 48.7014689167, 22.7097031285, -41.1402973647, -21.5570685361, -44.0503524604};
test_label[75] = '{48.7014689167};
test_output[75] = '{2.66564516973e-05};
############ END DEBUG ############*/
test_input[608:615] = '{32'hc2c25819, 32'hc216119b, 32'hc2b08f40, 32'hc259c585, 32'h42a994d7, 32'hc27a83cf, 32'h4212b0a5, 32'h4261cd2c};
test_label[76] = '{32'h4212b0a5};
test_output[76] = '{32'h42407909};
/*############ DEBUG ############
test_input[608:615] = '{-97.1720657879, -37.5171934029, -88.2797883787, -54.4428905929, 84.7907043818, -62.6287207806, 36.6725046033, 56.450362504};
test_label[76] = '{36.6725046033};
test_output[76] = '{48.1181997785};
############ END DEBUG ############*/
test_input[616:623] = '{32'hc1db0e8c, 32'h410eabfb, 32'hc12ce69c, 32'h414e51e8, 32'hc2b2587d, 32'hc280e0a0, 32'h41b6e37d, 32'h41c4ff07};
test_label[77] = '{32'hc2b2587d};
test_output[77] = '{32'h42e3e945};
/*############ DEBUG ############
test_input[616:623] = '{-27.3821024137, 8.91698706825, -10.8063012675, 12.8949969131, -89.1728263791, -64.4387218076, 22.8610784952, 24.6245255552};
test_label[77] = '{-89.1728263791};
test_output[77] = '{113.955603655};
############ END DEBUG ############*/
test_input[624:631] = '{32'hc25350d0, 32'hc28aa3ed, 32'hc0bb8fcf, 32'hc1fb316d, 32'h42a412cc, 32'hc2ba45d4, 32'hc21b8d88, 32'hc0c4e87f};
test_label[78] = '{32'hc25350d0};
test_output[78] = '{32'h4306dd9a};
/*############ DEBUG ############
test_input[624:631] = '{-52.8289191264, -69.3201666783, -5.86130474231, -31.3991331358, 82.036710407, -93.1363847315, -38.888214765, -6.15338103687};
test_label[78] = '{-52.8289191264};
test_output[78] = '{134.865629533};
############ END DEBUG ############*/
test_input[632:639] = '{32'h42235e0e, 32'h42b62e09, 32'hc2c7645a, 32'h4245d83a, 32'hc2789be6, 32'hc24205eb, 32'hc033ffae, 32'hc1ad7a21};
test_label[79] = '{32'hc1ad7a21};
test_output[79] = '{32'h42e18c91};
/*############ DEBUG ############
test_input[632:639] = '{40.8418519316, 91.0899113808, -99.6960011712, 49.4611593465, -62.1522443072, -48.5057777763, -2.81248036358, -21.6846327913};
test_label[79] = '{-21.6846327913};
test_output[79] = '{112.774544172};
############ END DEBUG ############*/
test_input[640:647] = '{32'h40d16ef6, 32'hc2c14e45, 32'hc21f7a9a, 32'hc28e3429, 32'h408305b8, 32'h40ebdd00, 32'h4141525c, 32'h423fd16d};
test_label[80] = '{32'hc21f7a9a};
test_output[80] = '{32'h42afa603};
/*############ DEBUG ############
test_input[640:647] = '{6.54479517708, -96.6528680396, -39.869726912, -71.1018722136, 4.09444812678, 7.37072749654, 12.0826076829, 47.9545180101};
test_label[80] = '{-39.869726912};
test_output[80] = '{87.8242449221};
############ END DEBUG ############*/
test_input[648:655] = '{32'h423cef1a, 32'h41e448b3, 32'hc20d32b3, 32'hc260e933, 32'hc1d13a04, 32'h42592766, 32'h42c1a1ee, 32'hc2c0130e};
test_label[81] = '{32'h42c1a1ee};
test_output[81] = '{32'h80000000};
/*############ DEBUG ############
test_input[648:655] = '{47.2334959802, 28.5354976169, -35.2995102595, -56.227732689, -26.153328143, 54.2884732716, 96.8162722323, -96.0372181639};
test_label[81] = '{96.8162722323};
test_output[81] = '{-0.0};
############ END DEBUG ############*/
test_input[656:663] = '{32'h4232ace0, 32'h4236c7fd, 32'hbfcbde48, 32'hc265f502, 32'hc1ee229c, 32'h42c31774, 32'hc28df0fc, 32'hc2bbfe5f};
test_label[82] = '{32'hbfcbde48};
test_output[82] = '{32'h42c646ed};
/*############ DEBUG ############
test_input[656:663] = '{44.6688232051, 45.6953021629, -1.59272097427, -57.4892670616, -29.7668993942, 97.5458036446, -70.9706731219, -93.9968167379};
test_label[82] = '{-1.59272097427};
test_output[82] = '{99.1385246189};
############ END DEBUG ############*/
test_input[664:671] = '{32'h425901bc, 32'hc13b7959, 32'hc2931f6d, 32'h42821081, 32'h428483ce, 32'h41efbbf4, 32'hc283cc2c, 32'h4229e117};
test_label[83] = '{32'h425901bc};
test_output[83] = '{32'h41443644};
/*############ DEBUG ############
test_input[664:671] = '{54.2516936806, -11.7171258548, -73.5613788818, 65.0322321451, 66.2574320671, 29.9667744011, -65.8987695416, 42.4698147483};
test_label[83] = '{54.2516936806};
test_output[83] = '{12.2632486484};
############ END DEBUG ############*/
test_input[672:679] = '{32'h4215fa92, 32'h42a65636, 32'hc2872e69, 32'h428584dc, 32'h429a5397, 32'hc16d6536, 32'h41a2bcd4, 32'h421ee818};
test_label[84] = '{32'h41a2bcd4};
test_output[84] = '{32'h427b5088};
/*############ DEBUG ############
test_input[672:679] = '{37.4946993383, 83.168382605, -67.5906457385, 66.7594901334, 77.1632587037, -14.8372098646, 20.3422017461, 39.7266557928};
test_label[84] = '{20.3422017461};
test_output[84] = '{62.8286439815};
############ END DEBUG ############*/
test_input[680:687] = '{32'hc2a30241, 32'h422e9382, 32'hc2276099, 32'h420fd334, 32'hc275af7c, 32'h428b3bfd, 32'hbf97c69f, 32'h42acde94};
test_label[85] = '{32'h420fd334};
test_output[85] = '{32'h4249e9f5};
/*############ DEBUG ############
test_input[680:687] = '{-81.5044018414, 43.6440514858, -41.8443318967, 35.9562531907, -61.4213724543, 69.6171629084, -1.18574891967, 86.434725863};
test_label[85] = '{35.9562531907};
test_output[85] = '{50.478472722};
############ END DEBUG ############*/
test_input[688:695] = '{32'h42949824, 32'h415d408d, 32'h42672579, 32'hc1bca46b, 32'h42aaea9b, 32'h41ad7ae4, 32'h41553104, 32'h42a3c9cd};
test_label[86] = '{32'h415d408d};
test_output[86] = '{32'h428f50d8};
/*############ DEBUG ############
test_input[688:695] = '{74.2971461744, 13.8282598291, 57.7865950301, -23.5802829736, 85.4582167651, 21.6850044935, 13.3244666641, 81.8941454121};
test_label[86] = '{13.8282598291};
test_output[86] = '{71.6579003494};
############ END DEBUG ############*/
test_input[696:703] = '{32'h422b153c, 32'h428ea8b0, 32'hc261b4e9, 32'h423608e8, 32'hc163890c, 32'hc143f41e, 32'hc2b60ff9, 32'h420dc47f};
test_label[87] = '{32'hc261b4e9};
test_output[87] = '{32'h42ff8324};
/*############ DEBUG ############
test_input[696:703] = '{42.7707350049, 71.3294640739, -56.4266703254, 45.5086957258, -14.2209587816, -12.247098643, -91.0311950736, 35.441890908};
test_label[87] = '{-56.4266703254};
test_output[87] = '{127.756134399};
############ END DEBUG ############*/
test_input[704:711] = '{32'h40928084, 32'hbeaa0fa7, 32'h4100fb5c, 32'h428ba456, 32'hc28d9aa5, 32'hc2b85d82, 32'h42c2a44a, 32'hc243d2be};
test_label[88] = '{32'hc2b85d82};
test_output[88] = '{32'h433d80e6};
/*############ DEBUG ############
test_input[704:711] = '{4.57818814785, -0.332150681874, 8.06136690952, 69.820969239, -70.8020383701, -92.1826320586, 97.3208742348, -48.9558039848};
test_label[88] = '{-92.1826320586};
test_output[88] = '{189.503506293};
############ END DEBUG ############*/
test_input[712:719] = '{32'hc2aaf83a, 32'h429e4570, 32'h42b78951, 32'hc1e3cb53, 32'h42001cb5, 32'hc2c6ba2d, 32'hc14b25d6, 32'h3fa149c3};
test_label[89] = '{32'hc2c6ba2d};
test_output[89] = '{32'h433f21bf};
/*############ DEBUG ############
test_input[712:719] = '{-85.4848191972, 79.1356212226, 91.7681930898, -28.4742796716, 32.0280325374, -99.3636276891, -12.6967371146, 1.26006352482};
test_label[89] = '{-99.3636276891};
test_output[89] = '{191.131824043};
############ END DEBUG ############*/
test_input[720:727] = '{32'hc243e11b, 32'h411b0c11, 32'hc2b4e6df, 32'h42377edf, 32'h42a7e3ce, 32'hc29a18be, 32'hc1394742, 32'h42632376};
test_label[90] = '{32'hc1394742};
test_output[90] = '{32'h42bf0cb7};
/*############ DEBUG ############
test_input[720:727] = '{-48.9698290958, 9.69044611786, -90.4509176428, 45.8738982777, 83.9449340964, -77.0483276363, -11.5798971906, 56.7846280428};
test_label[90] = '{-11.5798971906};
test_output[90] = '{95.524831287};
############ END DEBUG ############*/
test_input[728:735] = '{32'hc2a4cda7, 32'h42912a9c, 32'h42b79ff0, 32'h42b6007c, 32'hc1b1a30b, 32'hc05a7ba0, 32'h42c6c3b6, 32'h425cc42b};
test_label[91] = '{32'hc1b1a30b};
test_output[91] = '{32'h42f32cdb};
/*############ DEBUG ############
test_input[728:735] = '{-82.4016647572, 72.5832200347, 91.8123743017, 91.0009446888, -22.2046114572, -3.41379553626, 99.3822511274, 55.1915694252};
test_label[91] = '{-22.2046114572};
test_output[91] = '{121.587607174};
############ END DEBUG ############*/
test_input[736:743] = '{32'hc1bdb60a, 32'hc1f0f072, 32'hc28caef9, 32'hc15d62d6, 32'hc1f8dc26, 32'hc1cb0a88, 32'hc0c7438d, 32'h42981086};
test_label[92] = '{32'hc15d62d6};
test_output[92] = '{32'h42b3bce1};
/*############ DEBUG ############
test_input[736:743] = '{-23.7138865695, -30.1174057241, -70.3417433346, -13.8366295022, -31.1074949533, -25.3801413921, -6.22699606779, 76.0322738368};
test_label[92] = '{-13.8366295022};
test_output[92] = '{89.868903339};
############ END DEBUG ############*/
test_input[744:751] = '{32'hc29773b5, 32'h41e15439, 32'hc28eceed, 32'hc285305b, 32'h4266dd45, 32'hc246a121, 32'hc2b10a1b, 32'h42c287ef};
test_label[93] = '{32'hc28eceed};
test_output[93] = '{32'h4328ab6e};
/*############ DEBUG ############
test_input[744:751] = '{-75.7259900599, 28.1661251046, -71.4041517548, -66.5944417718, 57.7160833217, -49.657350664, -88.5197388478, 97.2654980071};
test_label[93] = '{-71.4041517548};
test_output[93] = '{168.669649762};
############ END DEBUG ############*/
test_input[752:759] = '{32'hc27e5377, 32'hc1306b7d, 32'hc27b92b6, 32'hc1ff1071, 32'hc206b374, 32'hc2329e16, 32'h4264f32c, 32'h41a3db78};
test_label[94] = '{32'hc206b374};
test_output[94] = '{32'h42b5d350};
/*############ DEBUG ############
test_input[752:759] = '{-63.5815081283, -11.0262421527, -62.8932737178, -31.883027111, -33.6752483334, -44.6543807391, 57.237472605, 20.4821624054};
test_label[94] = '{-33.6752483334};
test_output[94] = '{90.9127209384};
############ END DEBUG ############*/
test_input[760:767] = '{32'h42917fab, 32'h419f2c24, 32'h41b5a29c, 32'h428275a4, 32'hc1c2d236, 32'hc2079b12, 32'h40358250, 32'h420673e0};
test_label[95] = '{32'h42917fab};
test_output[95] = '{32'h3a0e2330};
/*############ DEBUG ############
test_input[760:767] = '{72.7493508928, 19.8965534911, 22.704400006, 65.2297673136, -24.3526420165, -33.9014345496, 2.83607872072, 33.6131572808};
test_label[95] = '{72.7493508928};
test_output[95] = '{0.000542211344978};
############ END DEBUG ############*/
test_input[768:775] = '{32'h421fa796, 32'hc16b465d, 32'hc1923058, 32'h4252a24b, 32'hc25fc5d7, 32'h41f83487, 32'hc2bdabb4, 32'hc1116ae3};
test_label[96] = '{32'hc1923058};
test_output[96] = '{32'h428ddd3c};
/*############ DEBUG ############
test_input[768:775] = '{39.9136589917, -14.7046788096, -18.2736052691, 52.6584899432, -55.9432036651, 31.0256477919, -94.8353587202, -9.08859577409};
test_label[96] = '{-18.2736052691};
test_output[96] = '{70.93209813};
############ END DEBUG ############*/
test_input[776:783] = '{32'h423ebb46, 32'hc2c23d26, 32'hc24e6f2c, 32'hc23c20e2, 32'hc1b447b8, 32'h41864f91, 32'hc1e074af, 32'h420b7b82};
test_label[97] = '{32'h41864f91};
test_output[97] = '{32'h41f726fd};
/*############ DEBUG ############
test_input[776:783] = '{47.6828854438, -97.119427991, -51.6085648792, -47.0321104701, -22.5350192936, 16.7888511643, -28.0569743408, 34.8706131881};
test_label[97] = '{16.7888511643};
test_output[97] = '{30.8940370066};
############ END DEBUG ############*/
test_input[784:791] = '{32'hc23c9721, 32'h42357999, 32'hc224f75f, 32'hc2030446, 32'h4251da66, 32'h42aa1b7c, 32'hc1bc719c, 32'h4197fc85};
test_label[98] = '{32'hc23c9721};
test_output[98] = '{32'h43043386};
/*############ DEBUG ############
test_input[784:791] = '{-47.1475877184, 45.3687461272, -41.2415748419, -32.7541738603, 52.4632788425, 85.0536784296, -23.5554731936, 18.9982997852};
test_label[98] = '{-47.1475877184};
test_output[98] = '{132.201266148};
############ END DEBUG ############*/
test_input[792:799] = '{32'h4239492a, 32'h4208d6fa, 32'hc2a23e2e, 32'hc2354b7c, 32'hc2c57813, 32'hc1acd49c, 32'hc264d94c, 32'hc23c8453};
test_label[99] = '{32'hc23c8453};
test_output[99] = '{32'h42bae6c0};
/*############ DEBUG ############
test_input[792:799] = '{46.3214496545, 34.2099387886, -81.121441623, -45.3237152104, -98.7345202138, -21.6038133378, -57.2122024064, -47.1292246996};
test_label[99] = '{-47.1292246996};
test_output[99] = '{93.4506798499};
############ END DEBUG ############*/
test_input[800:807] = '{32'h4251f069, 32'hc0391eb4, 32'hc28c8e55, 32'h413e3147, 32'hc1dc5717, 32'hc299da8d, 32'hc21cebfd, 32'h428b2b6e};
test_label[100] = '{32'hc0391eb4};
test_output[100] = '{32'h4290f463};
/*############ DEBUG ############
test_input[800:807] = '{52.4847741281, -2.89249906121, -70.2779920161, 11.8870305472, -27.5425236324, -76.9268533421, -39.2304583355, 69.5848214475};
test_label[100] = '{-2.89249906121};
test_output[100] = '{72.4773205461};
############ END DEBUG ############*/
test_input[808:815] = '{32'h419ccf4a, 32'hc2ae3bc8, 32'h429e44ac, 32'hc28cf24b, 32'hc2b0f2e2, 32'hc233e107, 32'hc214e4f9, 32'hc2aab339};
test_label[101] = '{32'hc214e4f9};
test_output[101] = '{32'h42e8b729};
/*############ DEBUG ############
test_input[808:815] = '{19.6012148534, -87.116760585, 79.1341265359, -70.4732321511, -88.4743828436, -44.9697542147, -37.2236063405, -85.3500454972};
test_label[101] = '{-37.2236063405};
test_output[101] = '{116.357732876};
############ END DEBUG ############*/
test_input[816:823] = '{32'h42a7fca1, 32'hc2831eb7, 32'hc2246506, 32'h42a118fe, 32'h416cc44b, 32'h421f9360, 32'h428eb999, 32'h41be7a9c};
test_label[102] = '{32'h42a7fca1};
test_output[102] = '{32'h3d00b422};
/*############ DEBUG ############
test_input[816:823] = '{83.993418133, -65.5599862537, -41.0986543934, 80.5488139533, 14.7979232095, 39.8939216235, 71.3624955838, 23.8098684372};
test_label[102] = '{83.993418133};
test_output[102] = '{0.0314217866164};
############ END DEBUG ############*/
test_input[824:831] = '{32'hc226453b, 32'h40e7b241, 32'hc282a089, 32'h427f26f8, 32'h425f8547, 32'h42bb2f6a, 32'hc227c142, 32'h3f275fb8};
test_label[103] = '{32'h40e7b241};
test_output[103] = '{32'h42acb446};
/*############ DEBUG ############
test_input[824:831] = '{-41.567609004, 7.24050970134, -65.3135469542, 63.788056545, 55.8801537271, 93.5926077146, -41.9387269286, 0.653804285052};
test_label[103] = '{7.24050970134};
test_output[103] = '{86.3520980132};
############ END DEBUG ############*/
test_input[832:839] = '{32'hc2c6cb3b, 32'h42840d6b, 32'h42372ffa, 32'hc18baed4, 32'hc283c64d, 32'hc169d876, 32'hc123aa1a, 32'h42b4170b};
test_label[104] = '{32'hc2c6cb3b};
test_output[104] = '{32'h433d7123};
/*############ DEBUG ############
test_input[832:839] = '{-99.3969351492, 66.0262091781, 45.7968535878, -17.4603655575, -65.8873075174, -14.6153465335, -10.2290289742, 90.0450058552};
test_label[104] = '{-99.3969351492};
test_output[104] = '{189.441941004};
############ END DEBUG ############*/
test_input[840:847] = '{32'hc2c6bbaa, 32'h4189f55d, 32'h41867ffb, 32'hc14fafe7, 32'h42aa4c3d, 32'h4163a623, 32'h429f02f0, 32'hc1617ef5};
test_label[105] = '{32'h429f02f0};
test_output[105] = '{32'h40b4b1bc};
/*############ DEBUG ############
test_input[840:847] = '{-99.3665281424, 17.2448061293, 16.8124899555, -12.980445028, 85.1489006694, 14.2280611133, 79.5057401583, -14.093495128};
test_label[105] = '{79.5057401583};
test_output[105] = '{5.64669591138};
############ END DEBUG ############*/
test_input[848:855] = '{32'hc2c368cd, 32'h42a9d717, 32'h4268f5d8, 32'h425573bf, 32'h42b77a5b, 32'hc2c21703, 32'h42aae042, 32'hc155715f};
test_label[106] = '{32'h42a9d717};
test_output[106] = '{32'h40da4c32};
/*############ DEBUG ############
test_input[848:855] = '{-97.7046903498, 84.9200990616, 58.2400829395, 53.3630338164, 91.7389769917, -97.0449460038, 85.4380004827, -13.3401781835};
test_label[106] = '{84.9200990616};
test_output[106] = '{6.82180111248};
############ END DEBUG ############*/
test_input[856:863] = '{32'hc292edce, 32'h40937978, 32'h42158604, 32'hc2bd19a4, 32'h42b768a7, 32'h42c1d369, 32'h42b11790, 32'h42961332};
test_label[107] = '{32'h42b768a7};
test_output[107] = '{32'h40a6dab4};
/*############ DEBUG ############
test_input[856:863] = '{-73.4644632701, 4.60857777063, 37.3808755224, -94.550078222, 91.7043989001, 96.9129101771, 88.5460200288, 75.0374898087};
test_label[107] = '{91.7043989001};
test_output[107] = '{5.21419732891};
############ END DEBUG ############*/
test_input[864:871] = '{32'hc1a2cce6, 32'hc1823432, 32'hc1383c90, 32'hc129e046, 32'hc25f043d, 32'hc2949b48, 32'hc2a090d9, 32'hc20a1b01};
test_label[108] = '{32'hc20a1b01};
test_output[108] = '{32'h41c2072d};
/*############ DEBUG ############
test_input[864:871] = '{-20.3500484098, -16.2754868886, -11.5147854329, -10.6172542615, -55.7541376452, -74.3032830463, -80.2829023838, -34.5263715797};
test_label[108] = '{-34.5263715797};
test_output[108] = '{24.2535029003};
############ END DEBUG ############*/
test_input[872:879] = '{32'hc2b46947, 32'hc24f237e, 32'hc04f5869, 32'h423a3495, 32'hc27f8b66, 32'h4258e243, 32'hc21e291f, 32'hc2aea02d};
test_label[109] = '{32'h4258e243};
test_output[109] = '{32'h39f4ae67};
/*############ DEBUG ############
test_input[872:879] = '{-90.2056164086, -51.7846591155, -3.23977113674, 46.551350192, -63.8861330934, 54.2209568597, -39.5401562079, -87.3128471125};
test_label[109] = '{54.2209568597};
test_output[109] = '{0.000466692477786};
############ END DEBUG ############*/
test_input[880:887] = '{32'hc2a65b84, 32'hc2051468, 32'hc2610173, 32'hc2b71185, 32'hc2bdec2f, 32'hc1d0c070, 32'h42bc2245, 32'hc2752d25};
test_label[110] = '{32'hc2bdec2f};
test_output[110] = '{32'h433d073a};
/*############ DEBUG ############
test_input[880:887] = '{-83.1787398367, -33.2699289323, -56.2514146174, -91.5342183263, -94.9612988389, -26.093963517, 94.0669296749, -61.2940871233};
test_label[110] = '{-94.9612988389};
test_output[110] = '{189.028228514};
############ END DEBUG ############*/
test_input[888:895] = '{32'hc297fadc, 32'h42a63671, 32'h4265a031, 32'h4186269e, 32'hc1c46809, 32'hc29ba37b, 32'hc2b58115, 32'h41133117};
test_label[111] = '{32'hc1c46809};
test_output[111] = '{32'h42d75073};
/*############ DEBUG ############
test_input[888:895] = '{-75.9899568427, 83.1063281479, 57.4064357101, 16.7688568567, -24.5507981468, -77.819293991, -90.7521126168, 9.19948485075};
test_label[111] = '{-24.5507981468};
test_output[111] = '{107.657126295};
############ END DEBUG ############*/
test_input[896:903] = '{32'h429a1bee, 32'hc288707e, 32'h42bf5f83, 32'hc2b87ee3, 32'h41c133a4, 32'hc1e56153, 32'h4274aeb1, 32'hc1e12730};
test_label[112] = '{32'hc2b87ee3};
test_output[112] = '{32'h433bef33};
/*############ DEBUG ############
test_input[896:903] = '{77.0545515039, -68.2197129191, 95.6865450838, -92.2478239877, 24.1502143507, -28.672522381, 61.1705961791, -28.1441346853};
test_label[112] = '{-92.2478239877};
test_output[112] = '{187.93436908};
############ END DEBUG ############*/
test_input[904:911] = '{32'h412f2d41, 32'hc274937f, 32'h42981cd7, 32'h42bd5fed, 32'hc25d3874, 32'hc1358dfd, 32'hc087dba6, 32'hc223ad15};
test_label[113] = '{32'hc1358dfd};
test_output[113] = '{32'h42d411ad};
/*############ DEBUG ############
test_input[904:911] = '{10.9485479612, -61.1440394247, 76.0563286029, 94.6873560786, -55.3051283037, -11.3471648979, -4.24556273823, -40.919027103};
test_label[113] = '{-11.3471648979};
test_output[113] = '{106.034520985};
############ END DEBUG ############*/
test_input[912:919] = '{32'h4191bfa2, 32'hc1f3d5b4, 32'hc2be4b19, 32'h42896b71, 32'hc14a9ade, 32'hc26e9532, 32'h4220e1e8, 32'h403fd006};
test_label[114] = '{32'hc2be4b19};
test_output[114] = '{32'h4323db45};
/*############ DEBUG ############
test_input[912:919] = '{18.2185709834, -30.4793468905, -95.1466784515, 68.7098466943, -12.6628094792, -59.6456999834, 40.2206120434, 2.99707171258};
test_label[114] = '{-95.1466784515};
test_output[114] = '{163.856525146};
############ END DEBUG ############*/
test_input[920:927] = '{32'hc23a0c01, 32'h42bd963a, 32'h41ba4e14, 32'h42c13061, 32'hbfa5765d, 32'hc020df49, 32'h42b8166f, 32'hc19c444b};
test_label[115] = '{32'h42b8166f};
test_output[115] = '{32'h4096ccfa};
/*############ DEBUG ############
test_input[920:927] = '{-46.5117226012, 94.7934119043, 23.2881246883, 96.5944925744, -1.29267462299, -2.5136283176, 92.0438178744, -19.5333468406};
test_label[115] = '{92.0438178744};
test_output[115] = '{4.71252176785};
############ END DEBUG ############*/
test_input[928:935] = '{32'hc2a179ca, 32'hc0e56925, 32'hc23c7ba7, 32'h41b81d15, 32'hc291e9a4, 32'h419a6c60, 32'h428892ee, 32'h424c5342};
test_label[116] = '{32'h41b81d15};
test_output[116] = '{32'h42351752};
/*############ DEBUG ############
test_input[928:935] = '{-80.7378706872, -7.16908518982, -47.1207532663, 23.0141998425, -72.9563259108, 19.3029174684, 68.286974392, 51.0813069468};
test_label[116] = '{23.0141998425};
test_output[116] = '{45.2727745832};
############ END DEBUG ############*/
test_input[936:943] = '{32'hc2b2cfb2, 32'h4239694f, 32'hc20adb6c, 32'h425b60fd, 32'h41c8dfe7, 32'hc290441c, 32'hc271e28d, 32'h42703c55};
test_label[117] = '{32'hc20adb6c};
test_output[117] = '{32'h42bd8ea8};
/*############ DEBUG ############
test_input[936:943] = '{-89.4056523174, 46.3528385869, -34.714280397, 54.8447152125, 25.1093275064, -72.1330237673, -60.471239476, 60.0589174553};
test_label[117] = '{-34.714280397};
test_output[117] = '{94.7786229958};
############ END DEBUG ############*/
test_input[944:951] = '{32'h410bf353, 32'h42c01a64, 32'h42c3d56c, 32'h42986b7e, 32'hc241e526, 32'h40ab5beb, 32'h42417def, 32'hc277ae55};
test_label[118] = '{32'h42417def};
test_output[118] = '{32'h4246c056};
/*############ DEBUG ############
test_input[944:951] = '{8.74690543358, 96.0515454476, 97.9168384319, 76.2099447382, -48.4737766184, 5.35497043263, 48.3729813385, -61.9202467184};
test_label[118] = '{48.3729813385};
test_output[118] = '{49.6878282816};
############ END DEBUG ############*/
test_input[952:959] = '{32'h42926ffc, 32'hc2b16926, 32'hc2697b42, 32'h41c14754, 32'h419dbbd3, 32'h42c10eab, 32'h41a3b322, 32'h3fcc440b};
test_label[119] = '{32'h41c14754};
test_output[119] = '{32'h4290bcd6};
/*############ DEBUG ############
test_input[952:959] = '{73.2187178089, -88.7053717703, -58.370367596, 24.1598286538, 19.7167117698, 96.5286509406, 20.4624678512, 1.59582655489};
test_label[119] = '{24.1598286538};
test_output[119] = '{72.3688222869};
############ END DEBUG ############*/
test_input[960:967] = '{32'h429f7f84, 32'h42846b07, 32'h4189b2d3, 32'h4286b74c, 32'hc2be2636, 32'h42250edf, 32'hc2a847c6, 32'h42bd1dbd};
test_label[120] = '{32'h42bd1dbd};
test_output[120] = '{32'h34c6c9c1};
/*############ DEBUG ############
test_input[960:967] = '{79.7490513499, 66.2090414843, 17.2123161423, 67.3580036932, -95.0746316331, 41.2645241294, -84.1401803227, 94.5580854438};
test_label[120] = '{94.5580854438};
test_output[120] = '{3.70271688915e-07};
############ END DEBUG ############*/
test_input[968:975] = '{32'h424941b1, 32'h420fa15e, 32'h4012453f, 32'h42b5ae9b, 32'hc29dcf78, 32'hc199fd2f, 32'h427c8b3f, 32'h4281b85d};
test_label[121] = '{32'h42b5ae9b};
test_output[121] = '{32'h2cd7e500};
/*############ DEBUG ############
test_input[968:975] = '{50.3141501107, 35.907583494, 2.28547653983, 90.8410265343, -78.9052115915, -19.2486253575, 63.1359832565, 64.8600869636};
test_label[121] = '{90.8410265343};
test_output[121] = '{6.13609163482e-12};
############ END DEBUG ############*/
test_input[976:983] = '{32'hc2890dd9, 32'hc1b953c0, 32'h424a597e, 32'hc0ed0f90, 32'hc297f72c, 32'hc2bdd6b0, 32'hc2873177, 32'hc1812baf};
test_label[122] = '{32'hc2bdd6b0};
test_output[122] = '{32'h431181b8};
/*############ DEBUG ############
test_input[976:983] = '{-68.5270488531, -23.1658928149, 50.5873929714, -7.40814953244, -75.9827600375, -94.9193142393, -67.596614524, -16.1463301691};
test_label[122] = '{-94.9193142393};
test_output[122] = '{145.506707211};
############ END DEBUG ############*/
test_input[984:991] = '{32'h429a242d, 32'hc28e38f5, 32'hc211b0a2, 32'hc02a9a06, 32'h41b7c5de, 32'h42ab5acd, 32'hc2af92b7, 32'hc2a26baa};
test_label[123] = '{32'hc2a26baa};
test_output[123] = '{32'h4326e347};
/*############ DEBUG ############
test_input[984:991] = '{77.0706576803, -71.1112444142, -36.4224913126, -2.66565076571, 22.9716146552, 85.6773449103, -87.7865544477, -81.2102799671};
test_label[123] = '{-81.2102799671};
test_output[123] = '{166.887807739};
############ END DEBUG ############*/
test_input[992:999] = '{32'hc242f21e, 32'hc1cdef32, 32'h4218930f, 32'hc264536a, 32'h41f9ac8f, 32'h42965b59, 32'hc202feb4, 32'hc2829b83};
test_label[124] = '{32'hc264536a};
test_output[124] = '{32'h43044287};
/*############ DEBUG ############
test_input[992:999] = '{-48.7364412998, -25.7417952206, 38.1436108392, -57.0814586463, 31.2092562036, 75.178412449, -32.748734587, -65.303735463};
test_label[124] = '{-57.0814586463};
test_output[124] = '{132.259871095};
############ END DEBUG ############*/
test_input[1000:1007] = '{32'h419f5e2a, 32'h42848b15, 32'hc2a17af3, 32'hc1bb2ce8, 32'h4184488f, 32'hc2820e69, 32'hc2c747d4, 32'h41630520};
test_label[125] = '{32'hc2820e69};
test_output[125] = '{32'h43034cbf};
/*############ DEBUG ############
test_input[1000:1007] = '{19.920977828, 66.2716478751, -80.7401359194, -23.3969272107, 16.5354297834, -65.0281478794, -99.6402925513, 14.188751127};
test_label[125] = '{-65.0281478794};
test_output[125] = '{131.299795754};
############ END DEBUG ############*/
test_input[1008:1015] = '{32'h4115eca9, 32'hc1c9f4c3, 32'hc1efa556, 32'hc124a7b1, 32'h41fdec42, 32'hc2c0a0bb, 32'hc29d27fa, 32'h42900491};
test_label[126] = '{32'hc29d27fa};
test_output[126] = '{32'h43169645};
/*############ DEBUG ############
test_input[1008:1015] = '{9.37027832693, -25.2445121218, -29.9557307414, -10.2909400718, 31.740360874, -96.3139261723, -78.5780793413, 72.0089165007};
test_label[126] = '{-78.5780793413};
test_output[126] = '{150.586995842};
############ END DEBUG ############*/
test_input[1016:1023] = '{32'h4293511f, 32'h42286435, 32'hc2928af7, 32'hc06263a4, 32'hbf8b3eb8, 32'h4295d70f, 32'h424cdcb6, 32'h42b494a0};
test_label[127] = '{32'h42b494a0};
test_output[127] = '{32'h349187ad};
/*############ DEBUG ############
test_input[1016:1023] = '{73.6584409758, 42.097859551, -73.2714171619, -3.53733155182, -1.08785157075, 74.9200361013, 51.2155398367, 90.2902805038};
test_label[127] = '{90.2902805038};
test_output[127] = '{2.71070722637e-07};
############ END DEBUG ############*/
test_input[1024:1031] = '{32'h4227a189, 32'hc1dbe710, 32'h412b929d, 32'hc29862cf, 32'hc1dc89c9, 32'h42a6d8b5, 32'hc2172eac, 32'h41ec5759};
test_label[128] = '{32'h41ec5759};
test_output[128] = '{32'h425785bd};
/*############ DEBUG ############
test_input[1024:1031] = '{41.9077481756, -27.4878241994, 10.7232944955, -76.1929854404, -27.5672770322, 83.4232563812, -37.7955772058, 29.5426509015};
test_label[128] = '{29.5426509015};
test_output[128] = '{53.8806054797};
############ END DEBUG ############*/
test_input[1032:1039] = '{32'hc27e9eb6, 32'hc2a92ce1, 32'hc2278b34, 32'hc2abad7a, 32'hc27a48c6, 32'hc2805832, 32'h422cee73, 32'h428da4ee};
test_label[129] = '{32'h422cee73};
test_output[129] = '{32'h41dcb6d2};
/*############ DEBUG ############
test_input[1032:1039] = '{-63.6549896308, -84.5876517632, -41.8859423758, -85.8388226929, -62.5710694409, -64.1722552563, 43.2328593718, 70.8221262214};
test_label[129] = '{43.2328593718};
test_output[129] = '{27.5892668497};
############ END DEBUG ############*/
test_input[1040:1047] = '{32'hc2649e63, 32'h415ed4fe, 32'hc299918b, 32'hc212a4ea, 32'hc263e23e, 32'hc216519a, 32'h418721a7, 32'hc061bc56};
test_label[130] = '{32'h418721a7};
test_output[130] = '{32'h3d4e0a9c};
/*############ DEBUG ############
test_input[1040:1047] = '{-57.1546747872, 13.9270001582, -76.7842651515, -36.6610499242, -56.9709377378, -37.579689629, 16.8914320728, -3.52712015775};
test_label[130] = '{16.8914320728};
test_output[130] = '{0.0503030854798};
############ END DEBUG ############*/
test_input[1048:1055] = '{32'h4235d12e, 32'h3ff94259, 32'h42849391, 32'h41e51d11, 32'hc28ab88e, 32'h42b05cd1, 32'hc2b311fc, 32'h3f0b1959};
test_label[131] = '{32'h42b05cd1};
test_output[131] = '{32'h2faaa8f4};
/*############ DEBUG ############
test_input[1048:1055] = '{45.4542753911, 1.94733729864, 66.2882124539, 28.6391924396, -69.3604561239, 88.181279451, -89.5351264198, 0.543355501518};
test_label[131] = '{88.181279451};
test_output[131] = '{3.10428682808e-10};
############ END DEBUG ############*/
test_input[1056:1063] = '{32'hc26b6de0, 32'h42913d6f, 32'hc1f77bd0, 32'hc288d019, 32'hc1f1d0d6, 32'hc2bed34a, 32'hc24eaf1b, 32'hc29c03b5};
test_label[132] = '{32'hc29c03b5};
test_output[132] = '{32'h4316a092};
/*############ DEBUG ############
test_input[1056:1063] = '{-58.8573002536, 72.6199837349, -30.9354555065, -68.4064392516, -30.226970269, -95.4126771244, -51.671001071, -78.0072414994};
test_label[132] = '{-78.0072414994};
test_output[132] = '{150.627225234};
############ END DEBUG ############*/
test_input[1064:1071] = '{32'h42223487, 32'hc273831a, 32'hc2801de8, 32'hc21673c1, 32'hc19e10fd, 32'hc292132f, 32'h42271d97, 32'h422c6e74};
test_label[133] = '{32'h42223487};
test_output[133] = '{32'h40367646};
/*############ DEBUG ############
test_input[1064:1071] = '{40.551295404, -60.8780285425, -64.0584133548, -37.6130403442, -19.7582950212, -73.0374676225, 41.7788953556, 43.1078642951};
test_label[133] = '{40.551295404};
test_output[133] = '{2.85096874684};
############ END DEBUG ############*/
test_input[1072:1079] = '{32'h41aaa51e, 32'hc24c3fc2, 32'h426002c8, 32'h42a3181a, 32'hc2862159, 32'h40577822, 32'hc101a10b, 32'hc198f798};
test_label[134] = '{32'h40577822};
test_output[134] = '{32'h429c5c59};
/*############ DEBUG ############
test_input[1072:1079] = '{21.3306230591, -51.062263719, 56.0027156578, 81.5470714502, -67.0651332863, 3.3667073973, -8.10181668772, -19.1208947066};
test_label[134] = '{3.3667073973};
test_output[134] = '{78.1803640529};
############ END DEBUG ############*/
test_input[1080:1087] = '{32'hc1515393, 32'h42c66549, 32'hc2a5cd52, 32'hc1b640c3, 32'h42c6d7ed, 32'hc252d5ee, 32'hc2459626, 32'h41f17f05};
test_label[135] = '{32'hc1515393};
test_output[135] = '{32'h42e22f25};
/*############ DEBUG ############
test_input[1080:1087] = '{-13.0829042562, 99.1978205816, -82.9010146626, -22.7816225268, 99.421732344, -52.7089167516, -49.396631121, 30.187020557};
test_label[135] = '{-13.0829042562};
test_output[135] = '{113.092081911};
############ END DEBUG ############*/
test_input[1088:1095] = '{32'hc2078443, 32'h41a45d96, 32'hc227960c, 32'hc2326278, 32'h42a58523, 32'h42addef1, 32'h413e3a72, 32'h42b647bc};
test_label[136] = '{32'h41a45d96};
test_output[136] = '{32'h428d380a};
/*############ DEBUG ############
test_input[1088:1095] = '{-33.8791617503, 20.5456961259, -41.8965306123, -44.5961616894, 82.7600305317, 86.9354321455, 11.8892687887, 91.1401074289};
test_label[136] = '{20.5456961259};
test_output[136] = '{70.6094526369};
############ END DEBUG ############*/
test_input[1096:1103] = '{32'hc20f8cf5, 32'hc2c1eac6, 32'h42664217, 32'hc2a98968, 32'hc223021b, 32'hc298d990, 32'h42c08420, 32'hc22847c7};
test_label[137] = '{32'hc2c1eac6};
test_output[137] = '{32'h43413773};
/*############ DEBUG ############
test_input[1096:1103] = '{-35.8876517533, -96.9585404576, 57.5645404363, -84.7683710492, -40.7520558592, -76.4249297013, 96.2580559804, -42.0700955342};
test_label[137] = '{-96.9585404576};
test_output[137] = '{193.216596438};
############ END DEBUG ############*/
test_input[1104:1111] = '{32'h41100fba, 32'hc2b2cd4c, 32'hc1e723a7, 32'hc2ab1235, 32'hc2a58823, 32'h42be38a0, 32'hc2653077, 32'h3e32b3df};
test_label[138] = '{32'hc2b2cd4c};
test_output[138] = '{32'h433882f6};
/*############ DEBUG ############
test_input[1104:1111] = '{9.00383981284, -89.4009736464, -28.8924078428, -85.5355612999, -82.7658912519, 95.1105964613, -57.2973287166, 0.174514284465};
test_label[138] = '{-89.4009736464};
test_output[138] = '{184.511570108};
############ END DEBUG ############*/
test_input[1112:1119] = '{32'h42159ed9, 32'h42ba9057, 32'hc270b9f2, 32'hc1b2b986, 32'h428480be, 32'hc2a8208b, 32'hc2597a56, 32'h42989376};
test_label[139] = '{32'hc1b2b986};
test_output[139] = '{32'h42e73eb9};
/*############ DEBUG ############
test_input[1112:1119] = '{37.4051260892, 93.281917188, -60.1815864055, -22.3405874964, 66.2514489265, -84.0635609765, -54.3694676297, 76.2880111892};
test_label[139] = '{-22.3405874964};
test_output[139] = '{115.622504726};
############ END DEBUG ############*/
test_input[1120:1127] = '{32'hc27dc130, 32'h405988d4, 32'h42b812fe, 32'h42ae0093, 32'hbf91430f, 32'h41fa738e, 32'hc2b0164b, 32'hc2ae262d};
test_label[140] = '{32'h41fa738e};
test_output[140] = '{32'h4272f2d8};
/*############ DEBUG ############
test_input[1120:1127] = '{-63.4386583091, 3.39897628355, 92.0370959369, 87.0011185665, -1.13485892154, 31.3064235478, -88.0435427362, -87.0745587279};
test_label[140] = '{31.3064235478};
test_output[140] = '{60.7371511984};
############ END DEBUG ############*/
test_input[1128:1135] = '{32'hc2874b83, 32'h427815c8, 32'h42ad94a5, 32'h41efb044, 32'hc2aaac6a, 32'hc1ec13b5, 32'hc20aac1e, 32'hc23024dd};
test_label[141] = '{32'h427815c8};
test_output[141] = '{32'h41c62703};
/*############ DEBUG ############
test_input[1128:1135] = '{-67.6474819073, 62.0212699595, 86.7903180131, 29.961067165, -85.3367497306, -29.5096220648, -34.6680831156, -44.0360000535};
test_label[141] = '{62.0212699595};
test_output[141] = '{24.7690480536};
############ END DEBUG ############*/
test_input[1136:1143] = '{32'h429c1105, 32'h41e80edf, 32'h429a477d, 32'hc203a719, 32'hc14385fa, 32'h41e23e64, 32'hc259b2a4, 32'h42a5dd06};
test_label[142] = '{32'h41e23e64};
test_output[142] = '{32'h425aa590};
/*############ DEBUG ############
test_input[1136:1143] = '{78.0332417426, 29.0072606236, 77.1396276311, -32.913182478, -12.2202087074, 28.2804634463, -54.4244540464, 82.931690046};
test_label[142] = '{28.2804634463};
test_output[142] = '{54.6616815841};
############ END DEBUG ############*/
test_input[1144:1151] = '{32'h42672d3e, 32'h428e037b, 32'hc23d821b, 32'hc25153b0, 32'h428a525a, 32'hc2232d21, 32'h42aa0b00, 32'hc266b7d3};
test_label[143] = '{32'hc25153b0};
test_output[143] = '{32'h43095a6c};
/*############ DEBUG ############
test_input[1144:1151] = '{57.7941825659, 71.0067959324, -47.3770550291, -52.3317275564, 69.1608394578, -40.7940706718, 85.0214858761, -57.6795173184};
test_label[143] = '{-52.3317275564};
test_output[143] = '{137.353214381};
############ END DEBUG ############*/
test_input[1152:1159] = '{32'h4285ccea, 32'hc2487609, 32'h4128bf72, 32'h416ed28e, 32'hc2709c7e, 32'hc239a624, 32'h42c28c32, 32'h42b5f90a};
test_label[144] = '{32'h4285ccea};
test_output[144] = '{32'h41f300f0};
/*############ DEBUG ############
test_input[1152:1159] = '{66.9002205626, -50.1152679106, 10.5467393441, 14.9264047814, -60.1528226155, -46.4122480367, 97.2738209136, 90.9864077435};
test_label[144] = '{66.9002205626};
test_output[144] = '{30.3754581882};
############ END DEBUG ############*/
test_input[1160:1167] = '{32'h42c3182e, 32'hc0845627, 32'hc23c362b, 32'h4207568d, 32'hc1d18cfb, 32'h401ba1d4, 32'hc273157d, 32'hc08dd63f};
test_label[145] = '{32'hc273157d};
test_output[145] = '{32'h431e5176};
/*############ DEBUG ############
test_input[1160:1167] = '{97.5472226303, -4.13551646818, -47.0528966476, 33.8345240745, -26.1938385965, 2.43175209068, -60.7709865288, -4.43240325912};
test_label[145] = '{-60.7709865288};
test_output[145] = '{158.318209159};
############ END DEBUG ############*/
test_input[1168:1175] = '{32'hc1d55b53, 32'hc0f3b40b, 32'hc2c78593, 32'hc299d4d2, 32'hc2898284, 32'hc2522550, 32'h42b6b046, 32'hc292eadc};
test_label[146] = '{32'hc2522550};
test_output[146] = '{32'h430fe177};
/*############ DEBUG ############
test_input[1168:1175] = '{-26.6695912574, -7.6157280076, -99.760887918, -76.9156669051, -68.7549145215, -52.5364381057, 91.3442828055, -73.458710623};
test_label[146] = '{-52.5364381057};
test_output[146] = '{143.880720911};
############ END DEBUG ############*/
test_input[1176:1183] = '{32'h421ff9bb, 32'hc2abf325, 32'h4281c35d, 32'hc27fa45e, 32'h4220d326, 32'h42c367f5, 32'hc19f4bdc, 32'hc2979214};
test_label[147] = '{32'hc2abf325};
test_output[147] = '{32'h4337ad8d};
/*############ DEBUG ############
test_input[1176:1183] = '{39.9938772035, -85.9748878915, 64.8815689925, -63.9105141298, 40.206199443, 97.7030396882, -19.9120414858, -75.7853107925};
test_label[147] = '{-85.9748878915};
test_output[147] = '{183.67792758};
############ END DEBUG ############*/
test_input[1184:1191] = '{32'hc2b45cdb, 32'h42933068, 32'hc2bf8189, 32'h4214a92a, 32'hc21e7652, 32'hc21533bb, 32'h416a4834, 32'h4294a9a0};
test_label[148] = '{32'hc2b45cdb};
test_output[148] = '{32'h4324e75f};
/*############ DEBUG ############
test_input[1184:1191] = '{-90.1813596891, 73.5945421914, -95.7530000771, 37.1652004452, -39.6155475048, -37.3005192535, 14.6426273696, 74.3312959389};
test_label[148] = '{-90.1813596891};
test_output[148] = '{164.903795461};
############ END DEBUG ############*/
test_input[1192:1199] = '{32'hc1cdb70e, 32'h42c3683f, 32'hc2c7fac6, 32'h422811ef, 32'hc14a2bb6, 32'h429e5a30, 32'h4200b911, 32'h414f0499};
test_label[149] = '{32'hc1cdb70e};
test_output[149] = '{32'h42f6d602};
/*############ DEBUG ############
test_input[1192:1199] = '{-25.7143821131, 97.7036051568, -99.9897931511, 42.0175131483, -12.6356718908, 79.1761471399, 32.180729137, 12.9386221094};
test_label[149] = '{-25.7143821131};
test_output[149] = '{123.417987279};
############ END DEBUG ############*/
test_input[1200:1207] = '{32'hc2333400, 32'h41aa7031, 32'hc28910a6, 32'hc1cf6619, 32'h4193bb22, 32'hc188a7a3, 32'hc1ec50ea, 32'h42bf54fc};
test_label[150] = '{32'hc1ec50ea};
test_output[150] = '{32'h42fa6937};
/*############ DEBUG ############
test_input[1200:1207] = '{-44.8007820002, 21.304780999, -68.5325127464, -25.9248523756, 18.466372978, -17.0818534385, -29.5395090268, 95.6659881264};
test_label[150] = '{-29.5395090268};
test_output[150] = '{125.205497153};
############ END DEBUG ############*/
test_input[1208:1215] = '{32'h42b8d37c, 32'h428d0484, 32'hc29cfde0, 32'hc1b0029b, 32'h41b966e5, 32'hc248d37e, 32'h429620c0, 32'h42860db9};
test_label[151] = '{32'hc29cfde0};
test_output[151] = '{32'h432ae8ae};
/*############ DEBUG ############
test_input[1208:1215] = '{92.413051997, 70.5088169369, -78.4958489032, -22.0012714632, 23.1752417827, -50.2065363816, 75.063965064, 67.0267994942};
test_label[151] = '{-78.4958489032};
test_output[151] = '{170.90890093};
############ END DEBUG ############*/
test_input[1216:1223] = '{32'hc16d0232, 32'h42b5ff6f, 32'hc28b5a87, 32'hc29756dc, 32'hc22200e3, 32'h42afd04d, 32'hc28d7cea, 32'hc19b14d0};
test_label[152] = '{32'hc19b14d0};
test_output[152] = '{32'h42dcdb5f};
/*############ DEBUG ############
test_input[1216:1223] = '{-14.8130363638, 90.9988914153, -69.6768076488, -75.669643992, -40.5008667781, 87.9068377466, -70.7439750001, -19.385161568};
test_label[152] = '{-19.385161568};
test_output[152] = '{110.428460801};
############ END DEBUG ############*/
test_input[1224:1231] = '{32'h4039d26f, 32'h41ea6227, 32'hc28a6d2a, 32'h41c7f99b, 32'hc2b8c0bf, 32'hc265d30b, 32'hc259251e, 32'h40ec6ea2};
test_label[153] = '{32'h41c7f99b};
test_output[153] = '{32'h408a107b};
/*############ DEBUG ############
test_input[1224:1231] = '{2.90346879846, 29.2979256973, -69.2132080638, 24.9968771541, -92.3764608099, -57.4560957841, -54.286247007, 7.38850521594};
test_label[153] = '{24.9968771541};
test_output[153] = '{4.31451184435};
############ END DEBUG ############*/
test_input[1232:1239] = '{32'h4168e937, 32'h42b79933, 32'hc229a093, 32'h42013fdf, 32'h412a1bed, 32'h41c7b28d, 32'h428482af, 32'h4284d2d4};
test_label[154] = '{32'h412a1bed};
test_output[154] = '{32'h42a255b5};
/*############ DEBUG ############
test_input[1232:1239] = '{14.5569372226, 91.799218374, -42.4068108369, 32.3123735205, 10.6318180535, 24.9621820698, 66.2552392298, 66.4117705991};
test_label[154] = '{10.6318180535};
test_output[154] = '{81.1674003204};
############ END DEBUG ############*/
test_input[1240:1247] = '{32'hc2c31d40, 32'hc289fcdb, 32'hc27ab0fd, 32'h41bdcd89, 32'h424689fd, 32'h42b42c74, 32'h4226f7b4, 32'hc281c554};
test_label[155] = '{32'hc281c554};
test_output[155] = '{32'h431af8e4};
/*############ DEBUG ############
test_input[1240:1247] = '{-97.5571322767, -68.9938587554, -62.6728389705, 23.7253593584, 49.634752655, 90.0868256246, 41.741898318, -64.8854084399};
test_label[155] = '{-64.8854084399};
test_output[155] = '{154.972234065};
############ END DEBUG ############*/
test_input[1248:1255] = '{32'h42c1db70, 32'h42bb1399, 32'h42417637, 32'h42a426ba, 32'hc15119aa, 32'hc2810ec5, 32'hc293361a, 32'hc1a59d0c};
test_label[156] = '{32'hc1a59d0c};
test_output[156] = '{32'h42eb53ab};
/*############ DEBUG ############
test_input[1248:1255] = '{96.9285924079, 93.5382745972, 48.3654457993, 82.0756405869, -13.0687660946, -64.5288445062, -73.605664667, -20.7016821563};
test_label[156] = '{-20.7016821563};
test_output[156] = '{117.663417538};
############ END DEBUG ############*/
test_input[1256:1263] = '{32'hc2b97a9f, 32'h4282e56e, 32'hc2a3ce08, 32'h414063a6, 32'h412d79cb, 32'hc23a31d3, 32'hc278ce83, 32'h411f9516};
test_label[157] = '{32'h412d79cb};
test_output[157] = '{32'h425a6c69};
/*############ DEBUG ############
test_input[1256:1263] = '{-92.7394940077, 65.4481028779, -81.9024042079, 12.0243277731, 10.84223459, -46.5486574232, -62.2016734841, 9.97389786617};
test_label[157] = '{10.84223459};
test_output[157] = '{54.6058682879};
############ END DEBUG ############*/
test_input[1264:1271] = '{32'h42788f93, 32'h42b7424f, 32'h42af4b8a, 32'h4287ddac, 32'hc29bafb4, 32'h429a54f6, 32'h41b21bd2, 32'h426a26f3};
test_label[158] = '{32'h42b7424f};
test_output[158] = '{32'h3c975e39};
/*############ DEBUG ############
test_input[1264:1271] = '{62.1402095396, 91.6295123139, 87.6475382718, 67.9329553422, -77.8431682161, 77.1659413605, 22.2635843385, 58.5380377606};
test_label[158] = '{91.6295123139};
test_output[158] = '{0.0184775464244};
############ END DEBUG ############*/
test_input[1272:1279] = '{32'h42784ca8, 32'h417b48e5, 32'hbf3112e8, 32'hc208bdea, 32'h4227dae3, 32'h424f9060, 32'hc2944b64, 32'h42af68b1};
test_label[159] = '{32'hc2944b64};
test_output[159] = '{32'h4321da0a};
/*############ DEBUG ############
test_input[1272:1279] = '{62.0748611893, 15.7052964963, -0.691694745524, -34.1854643196, 41.9637558265, 51.8909899717, -74.1472461227, 87.7044735603};
test_label[159] = '{-74.1472461227};
test_output[159] = '{161.851719683};
############ END DEBUG ############*/
test_input[1280:1287] = '{32'h410fa503, 32'hc2423e23, 32'h429b47b2, 32'hc2b05ee1, 32'h41cd350a, 32'hc11ec9d2, 32'h425a17ce, 32'hc2311be7};
test_label[160] = '{32'hc2b05ee1};
test_output[160] = '{32'h4325d34a};
/*############ DEBUG ############
test_input[1280:1287] = '{8.97778641697, -48.5606804234, 77.6400336381, -88.1853117152, 25.6508983272, -9.9242723372, 54.5232463919, -44.2772502844};
test_label[160] = '{-88.1853117152};
test_output[160] = '{165.825345353};
############ END DEBUG ############*/
test_input[1288:1295] = '{32'hbe976d47, 32'h420ab26f, 32'h42b65ac2, 32'h41614a71, 32'h428a304f, 32'hc29f4b24, 32'h4113398f, 32'h41e4ffb2};
test_label[161] = '{32'h4113398f};
test_output[161] = '{32'h42a3f390};
/*############ DEBUG ############
test_input[1288:1295] = '{-0.295755593215, 34.674251512, 91.1772637598, 14.0806744508, 69.0943558515, -79.6467626459, 9.20155198877, 28.6248506744};
test_label[161] = '{9.20155198877};
test_output[161] = '{81.9757117713};
############ END DEBUG ############*/
test_input[1296:1303] = '{32'h428cf4e6, 32'hc2a4e279, 32'hc1b3f4b6, 32'h42a3cae7, 32'h42aadfda, 32'hc29ae8e3, 32'h424fb4c5, 32'hc285eb89};
test_label[162] = '{32'h428cf4e6};
test_output[162] = '{32'h416fccab};
/*############ DEBUG ############
test_input[1296:1303] = '{70.4783173403, -82.4423257838, -22.4944876615, 81.8962939712, 85.4372101407, -77.4548557822, 51.9265321152, -66.9600298428};
test_label[162] = '{70.4783173403};
test_output[162] = '{14.9874676983};
############ END DEBUG ############*/
test_input[1304:1311] = '{32'h41e407fe, 32'hc294cf01, 32'hc18ec3e8, 32'hc29dda35, 32'h422b3387, 32'hbfefbc5f, 32'hc2310dc9, 32'hc281ced4};
test_label[163] = '{32'hc2310dc9};
test_output[163] = '{32'h42ae20a8};
/*############ DEBUG ############
test_input[1304:1311] = '{28.5039023734, -74.4043009361, -17.8456582698, -78.9261869586, 42.8003189424, -1.87293611376, -44.2634638083, -64.9039610899};
test_label[163] = '{-44.2634638083};
test_output[163] = '{87.0637833689};
############ END DEBUG ############*/
test_input[1312:1319] = '{32'hc233e50f, 32'hc22ebd49, 32'hc231df24, 32'h41d28023, 32'hc18ab9cc, 32'hc1ea7e08, 32'h4202554a, 32'hc22a327c};
test_label[164] = '{32'h41d28023};
test_output[164] = '{32'h40c8b93c};
/*############ DEBUG ############
test_input[1312:1319] = '{-44.9736889793, -43.6848486812, -44.4679103266, 26.3125670889, -17.3407218266, -29.3115384531, 32.5832898662, -42.5493006775};
test_label[164] = '{26.3125670889};
test_output[164] = '{6.2726118533};
############ END DEBUG ############*/
test_input[1320:1327] = '{32'h42af8b5c, 32'hc23c7065, 32'h423f518d, 32'hc29177e2, 32'hc21bd825, 32'hc1a6d1bf, 32'h4251607a, 32'h42b6508a};
test_label[165] = '{32'h423f518d};
test_output[165] = '{32'h422d71a4};
/*############ DEBUG ############
test_input[1320:1327] = '{87.7721840118, -47.1097597517, 47.8296383867, -72.7341443739, -38.9610804029, -20.8524152341, 52.344215906, 91.157302827};
test_label[165] = '{47.8296383867};
test_output[165] = '{43.360976982};
############ END DEBUG ############*/
test_input[1328:1335] = '{32'h426d3009, 32'hc25b299d, 32'h423dcaa2, 32'h428f5db6, 32'h41d2bd44, 32'h3f4febbf, 32'hc2294bd3, 32'h42bdb313};
test_label[166] = '{32'h42bdb313};
test_output[166] = '{32'h2ebf0200};
/*############ DEBUG ############
test_input[1328:1335] = '{59.2969077446, -54.7906385834, 47.4478847107, 71.6830302089, 26.3424144577, 0.812190951027, -42.3240482521, 94.8497547254};
test_label[166] = '{94.8497547254};
test_output[166] = '{8.68602967368e-11};
############ END DEBUG ############*/
test_input[1336:1343] = '{32'h418f294c, 32'hc0d3f356, 32'hc291bf87, 32'hc2933ef8, 32'hc2c0b115, 32'hc2573d41, 32'h41ef7213, 32'h4226f117};
test_label[167] = '{32'h41ef7213};
test_output[167] = '{32'h413ce03e};
/*############ DEBUG ############
test_input[1336:1343] = '{17.895163828, -6.62345389313, -72.8740750521, -73.6229859122, -96.3458634015, -53.8098190123, 29.9307002806, 41.7354395209};
test_label[167] = '{29.9307002806};
test_output[167] = '{11.8047467094};
############ END DEBUG ############*/
test_input[1344:1351] = '{32'hbda29ab0, 32'h40dee5fe, 32'h429a807e, 32'hc2832cfb, 32'h42126814, 32'hc1ee386b, 32'hc228e423, 32'hc29e19a0};
test_label[168] = '{32'hc2832cfb};
test_output[168] = '{32'h430ed6bc};
/*############ DEBUG ############
test_input[1344:1351] = '{-0.0793966019769, 6.96557519478, 77.2509605163, -65.5878527826, 36.6016389104, -29.7775476401, -42.2227892201, -79.0500471052};
test_label[168] = '{-65.5878527826};
test_output[168] = '{142.838813299};
############ END DEBUG ############*/
test_input[1352:1359] = '{32'h4121a165, 32'hc250c25e, 32'h41f55c76, 32'h422a0ba0, 32'h42acb850, 32'h4298b598, 32'hc182ea9c, 32'h402e5480};
test_label[169] = '{32'h4298b598};
test_output[169] = '{32'h412015ef};
/*############ DEBUG ############
test_input[1352:1359] = '{10.101902963, -52.1898121885, 30.6701472805, 42.51135177, 86.3599880312, 76.354678612, -16.3645558957, 2.72390753958};
test_label[169] = '{76.354678612};
test_output[169] = '{10.0053545777};
############ END DEBUG ############*/
test_input[1360:1367] = '{32'h425a21f8, 32'hc28ba3d0, 32'hc1f4ad80, 32'h41df957d, 32'hc01aa6c1, 32'h4226b6e5, 32'h41beaec0, 32'hc262e1d3};
test_label[170] = '{32'h4226b6e5};
test_output[170] = '{32'h414dac4f};
/*############ DEBUG ############
test_input[1360:1367] = '{54.5331723119, -69.8199460544, -30.5847169907, 27.9479924736, -2.41642777916, 41.6786075448, 23.8353273544, -56.7205331584};
test_label[170] = '{41.6786075448};
test_output[170] = '{12.8545673812};
############ END DEBUG ############*/
test_input[1368:1375] = '{32'hc0e89c88, 32'h41862f44, 32'hbfd3fdc7, 32'hc29a9bf2, 32'h42c323fb, 32'hc1c6d02c, 32'hc1d49e54, 32'h413c397b};
test_label[171] = '{32'h42c323fb};
test_output[171] = '{32'h80000000};
/*############ DEBUG ############
test_input[1368:1375] = '{-7.26910791047, 16.7730798647, -1.65618213495, -77.3045842043, 97.5702762848, -24.8516473339, -26.5773086939, 11.7640330274};
test_label[171] = '{97.5702762848};
test_output[171] = '{-0.0};
############ END DEBUG ############*/
test_input[1376:1383] = '{32'hc207bdaa, 32'h4239b399, 32'h42387f66, 32'h423fe2bd, 32'hc1903d81, 32'hc2be37c8, 32'h4239ea1a, 32'hc2b89626};
test_label[172] = '{32'h423fe2bd};
test_output[172] = '{32'h3eef3663};
/*############ DEBUG ############
test_input[1376:1383] = '{-33.9352179867, 46.425390225, 46.1244116522, 47.9714238998, -18.0300320983, -95.1089487691, 46.4786136263, -92.2932551407};
test_label[172] = '{47.9714238998};
test_output[172] = '{0.467211817273};
############ END DEBUG ############*/
test_input[1384:1391] = '{32'h421f5a27, 32'hc180bda0, 32'hc28fbfd1, 32'h41cacad9, 32'hc0dbe018, 32'h42c09ae8, 32'h42b90921, 32'hc2612b5d};
test_label[173] = '{32'hc2612b5d};
test_output[173] = '{32'h43189e0b};
/*############ DEBUG ############
test_input[1384:1391] = '{39.8380385838, -16.0925909416, -71.8746399678, 25.3490472847, -6.87110499816, 96.3025487298, 92.5178335134, -56.2923466981};
test_label[173] = '{-56.2923466981};
test_output[173] = '{152.617356607};
############ END DEBUG ############*/
test_input[1392:1399] = '{32'h42a1ae6f, 32'hc2c5b87a, 32'h420616e2, 32'hc29a66d5, 32'hc14e6716, 32'h428f9dce, 32'hc1efaa8c, 32'h425157f4};
test_label[174] = '{32'hc14e6716};
test_output[174] = '{32'h42bb7b61};
/*############ DEBUG ############
test_input[1392:1399] = '{80.8406908886, -98.8603066354, 33.5223480706, -77.2008443623, -12.9001672509, 71.8082111003, -29.9582755657, 52.3358920488};
test_label[174] = '{-12.9001672509};
test_output[174] = '{93.7409775983};
############ END DEBUG ############*/
test_input[1400:1407] = '{32'hc2a61d44, 32'h42a54a38, 32'h42aeb3cf, 32'hc2aedd9c, 32'h42bf60ff, 32'hc1a99b42, 32'h41cb6bb2, 32'h427b5746};
test_label[175] = '{32'hc2aedd9c};
test_output[175] = '{32'h43371f5d};
/*############ DEBUG ############
test_input[1400:1407] = '{-83.0571592236, 82.6449560268, 87.3511870405, -87.4328282203, 95.6894467311, -21.2008086668, 25.4275860086, 62.8352264609};
test_label[175] = '{-87.4328282203};
test_output[175] = '{183.122516272};
############ END DEBUG ############*/
test_input[1408:1415] = '{32'h424f324c, 32'h41f8d0fd, 32'h42b30b68, 32'h42c57b0c, 32'hc2aaf22c, 32'h429ba21e, 32'h42b6e756, 32'h41d6a518};
test_label[176] = '{32'h424f324c};
test_output[176] = '{32'h423bc49a};
/*############ DEBUG ############
test_input[1408:1415] = '{51.7991172471, 31.1020458297, 89.5222747329, 98.7403281709, -85.472995352, 77.8166325155, 91.4518296966, 26.8306124063};
test_label[176] = '{51.7991172471};
test_output[176] = '{46.9419932035};
############ END DEBUG ############*/
test_input[1416:1423] = '{32'hc2858e32, 32'hc1a1b9fc, 32'h429429e1, 32'h42c7a9a1, 32'hc275687f, 32'h4171e9be, 32'h41d64607, 32'h42b57825};
test_label[177] = '{32'hc2858e32};
test_output[177] = '{32'h43269bf1};
/*############ DEBUG ############
test_input[1416:1423] = '{-66.7777282573, -20.2158131053, 74.0817916919, 99.8313098593, -61.3520461255, 15.1195657746, 26.784193829, 90.7346542949};
test_label[177] = '{-66.7777282573};
test_output[177] = '{166.60915015};
############ END DEBUG ############*/
test_input[1424:1431] = '{32'hc2bc7dbd, 32'h428fd054, 32'h4282a0ae, 32'hc286c26c, 32'h41bac100, 32'hc1f43608, 32'h41312a37, 32'hc0978938};
test_label[178] = '{32'hc0978938};
test_output[178] = '{32'h4299499b};
/*############ DEBUG ############
test_input[1424:1431] = '{-94.2455846059, 71.9068931771, 65.3138255494, -67.379729847, 23.3442380443, -30.5263825499, 11.0728067821, -4.73550038721};
test_label[178] = '{-4.73550038721};
test_output[178] = '{76.6437624583};
############ END DEBUG ############*/
test_input[1432:1439] = '{32'hc18b89c9, 32'h429e27e6, 32'hc29eb4c7, 32'h41b9f508, 32'h41e6a621, 32'h42b117cc, 32'hc0f48a40, 32'hc2b3eeb0};
test_label[179] = '{32'h42b117cc};
test_output[179] = '{32'h38a1fbbf};
/*############ DEBUG ############
test_input[1432:1439] = '{-17.442277824, 79.0779233974, -79.35308187, 23.2446445631, 28.8311175195, 88.5464818426, -7.64187634024, -89.9661849541};
test_label[179] = '{88.5464818426};
test_output[179] = '{7.7239693754e-05};
############ END DEBUG ############*/
test_input[1440:1447] = '{32'hc1afb708, 32'h42a404f5, 32'hc29341d6, 32'hc27f8d1e, 32'h426fe63a, 32'hc2b38795, 32'hc281f8f5, 32'hc2a261c1};
test_label[180] = '{32'hc29341d6};
test_output[180] = '{32'h431ba366};
/*############ DEBUG ############
test_input[1440:1447] = '{-21.9643709778, 82.0096828029, -73.6285861839, -63.8878106247, 59.9748294857, -89.7648082972, -64.9862441053, -81.1909262902};
test_label[180] = '{-73.6285861839};
test_output[180] = '{155.638268987};
############ END DEBUG ############*/
test_input[1448:1455] = '{32'h42a29568, 32'hc005d3d9, 32'h41cfa6ec, 32'hc14c22db, 32'hc2b45951, 32'h4241b024, 32'h41ad107a, 32'hc22a88aa};
test_label[181] = '{32'hc22a88aa};
test_output[181] = '{32'h42f7d9bd};
/*############ DEBUG ############
test_input[1448:1455] = '{81.291811867, -2.09105508451, 25.9565057632, -12.7585094792, -90.174447423, 48.4220127103, 21.6330444335, -42.6334592262};
test_label[181] = '{-42.6334592262};
test_output[181] = '{123.925271093};
############ END DEBUG ############*/
test_input[1456:1463] = '{32'hc26c4716, 32'hc29619cb, 32'h42939fb5, 32'hc2439ce7, 32'hc1b6151e, 32'h42a2d6fa, 32'hc1876db1, 32'hc1eb141c};
test_label[182] = '{32'h42939fb5};
test_output[182] = '{32'h40f37863};
/*############ DEBUG ############
test_input[1456:1463] = '{-59.0694189765, -75.050377975, 73.8119303249, -48.903224797, -22.7603103685, 81.4198796487, -16.9285595974, -29.3848195294};
test_label[182] = '{73.8119303249};
test_output[182] = '{7.60844568958};
############ END DEBUG ############*/
test_input[1464:1471] = '{32'h41c65e7a, 32'hc298c9e1, 32'hc1b3f544, 32'hc11028fd, 32'hc249d85f, 32'h42373ca1, 32'h4274182e, 32'h419e7a04};
test_label[183] = '{32'hc298c9e1};
test_output[183] = '{32'h43096afc};
/*############ DEBUG ############
test_input[1464:1471] = '{24.7961302461, -76.3942952055, -22.4947580815, -9.01000662646, -50.4612995923, 45.8092072453, 61.02361355, 19.8095773749};
test_label[183] = '{-76.3942952055};
test_output[183] = '{137.417909002};
############ END DEBUG ############*/
test_input[1472:1479] = '{32'hc28170b2, 32'hc18ecf86, 32'hc28e5e96, 32'hc1d0138d, 32'h429e3808, 32'hc2208f7a, 32'h427f59fc, 32'hc23e7d02};
test_label[184] = '{32'h429e3808};
test_output[184] = '{32'h347a595f};
/*############ DEBUG ############
test_input[1472:1479] = '{-64.7201097659, -17.8513295657, -71.1847408139, -26.0095461612, 79.109434359, -40.1401151929, 63.8378754417, -47.6220783362};
test_label[184] = '{79.109434359};
test_output[184] = '{2.33155777443e-07};
############ END DEBUG ############*/
test_input[1480:1487] = '{32'hc1f7929f, 32'hc2920cd0, 32'h42b4c74e, 32'hc27a80e1, 32'hc29109a5, 32'hc1b3cce0, 32'h41ba60c9, 32'h42c5b771};
test_label[185] = '{32'hc1b3cce0};
test_output[185] = '{32'h42f2aac4};
/*############ DEBUG ############
test_input[1480:1487] = '{-30.9465919454, -73.0250282189, 90.3892643527, -62.6258601116, -72.5188333048, -22.4750365509, 23.2972580128, 98.8582806103};
test_label[185] = '{-22.4750365509};
test_output[185] = '{121.33352701};
############ END DEBUG ############*/
test_input[1488:1495] = '{32'hc2a01dc7, 32'hc1cb6a41, 32'hc2898efe, 32'hc291e97b, 32'h42ab343a, 32'h41815428, 32'hc1d33151, 32'hc2b8fa52};
test_label[186] = '{32'hc291e97b};
test_output[186] = '{32'h431e8eda};
/*############ DEBUG ############
test_input[1488:1495] = '{-80.0581604573, -25.4268823882, -68.7792807574, -72.9560164637, 85.6020022689, 16.1660928178, -26.3990800939, -92.4889055362};
test_label[186] = '{-72.9560164637};
test_output[186] = '{158.558018733};
############ END DEBUG ############*/
test_input[1496:1503] = '{32'hc293d8f4, 32'hc28cb1cb, 32'h413b634e, 32'h42b7fc28, 32'hc2b60d7e, 32'h421ea5f7, 32'h42321227, 32'hc2359607};
test_label[187] = '{32'h421ea5f7};
test_output[187] = '{32'h42515258};
/*############ DEBUG ############
test_input[1496:1503] = '{-73.9237368494, -70.347249796, 11.7117443673, 91.992491064, -91.0263545429, 39.6620767039, 44.517725142, -45.3965103253};
test_label[187] = '{39.6620767039};
test_output[187] = '{52.3304143602};
############ END DEBUG ############*/
test_input[1504:1511] = '{32'h42af55c4, 32'hc112098e, 32'hc1a92148, 32'hc2735b3d, 32'hc2764f4c, 32'hc292f486, 32'hc1b2542c, 32'hc2a508f6};
test_label[188] = '{32'hc2735b3d};
test_output[188] = '{32'h431481b1};
/*############ DEBUG ############
test_input[1504:1511] = '{87.6675077362, -9.12733251096, -21.1412503542, -60.8390993607, -61.5774389312, -73.4775815295, -22.2910988685, -82.5175035516};
test_label[188] = '{-60.8390993607};
test_output[188] = '{148.506607097};
############ END DEBUG ############*/
test_input[1512:1519] = '{32'h42815f8d, 32'hc0ff65d2, 32'hc2b80968, 32'hc248b194, 32'hc19e656a, 32'h4200ccff, 32'hc2896df4, 32'hc2c6dbfa};
test_label[189] = '{32'hc2896df4};
test_output[189] = '{32'h430566c1};
/*############ DEBUG ############
test_input[1512:1519] = '{64.6866247466, -7.98117928046, -92.0183713942, -50.173415529, -19.7995194193, 32.2001930777, -68.7147545582, -99.4296426581};
test_label[189] = '{-68.7147545582};
test_output[189] = '{133.401379305};
############ END DEBUG ############*/
test_input[1520:1527] = '{32'h429dcbf2, 32'hc234b6fa, 32'hc22acccf, 32'hc2b82ff9, 32'hc1b7dc62, 32'h41f19cac, 32'hc28fbad4, 32'h42c19d04};
test_label[190] = '{32'h429dcbf2};
test_output[190] = '{32'h418f4449};
/*############ DEBUG ############
test_input[1520:1527] = '{78.8983271302, -45.1786898897, -42.7000102265, -92.0936938791, -22.9826093171, 30.2014999566, -71.864901346, 96.8066691426};
test_label[190] = '{78.8983271302};
test_output[190] = '{17.9083420291};
############ END DEBUG ############*/
test_input[1528:1535] = '{32'h41a23a8d, 32'hc261c41c, 32'hc2a22087, 32'hc2996b70, 32'hc19ce51c, 32'h42b2681e, 32'h42942eb3, 32'h41b77c5d};
test_label[191] = '{32'hc19ce51c};
test_output[191] = '{32'h42d9a165};
/*############ DEBUG ############
test_input[1528:1535] = '{20.2785900037, -56.4415131856, -81.0635273269, -76.7098355582, -19.6118694747, 89.2033542864, 74.0912103941, 22.9357246458};
test_label[191] = '{-19.6118694747};
test_output[191] = '{108.815224035};
############ END DEBUG ############*/
test_input[1536:1543] = '{32'hc14cd827, 32'h42342a40, 32'h4291c9bb, 32'hc1bbac7d, 32'hc2314080, 32'h422292b3, 32'hc2a4e45c, 32'h4174848f};
test_label[192] = '{32'h422292b3};
test_output[192] = '{32'h420100c3};
/*############ DEBUG ############
test_input[1536:1543] = '{-12.8027713066, 45.0412584773, 72.8940028631, -23.4592226723, -44.3129901542, 40.6432592733, -82.4460152849, 15.2823633685};
test_label[192] = '{40.6432592733};
test_output[192] = '{32.2507435898};
############ END DEBUG ############*/
test_input[1544:1551] = '{32'hc29b4bc9, 32'h424b9b61, 32'h42aab031, 32'h428a3000, 32'h42b6aded, 32'h4278471a, 32'hc16784f7, 32'hc2453ed5};
test_label[193] = '{32'hc2453ed5};
test_output[193] = '{32'h430ca74f};
/*############ DEBUG ############
test_input[1544:1551] = '{-77.6480209634, 50.9017360208, 85.3441270565, 69.0937516066, 91.3396999623, 62.06943548, -14.4699625569, -49.3113602679};
test_label[193] = '{-49.3113602679};
test_output[193] = '{140.653546886};
############ END DEBUG ############*/
test_input[1552:1559] = '{32'hc25bd824, 32'h41df36d6, 32'h4272dc49, 32'hc1d42176, 32'hc2addeaf, 32'h42b38d3d, 32'h42982ddb, 32'h4259ef72};
test_label[194] = '{32'h42b38d3d};
test_output[194] = '{32'h3598bb0e};
/*############ DEBUG ############
test_input[1552:1559] = '{-54.9610764383, 27.9017759032, 60.7151208393, -26.5163377363, -86.934925115, 89.7758560097, 76.0895586192, 54.4838333943};
test_label[194] = '{89.7758560097};
test_output[194] = '{1.13793226094e-06};
############ END DEBUG ############*/
test_input[1560:1567] = '{32'hc29b15fb, 32'h410b806e, 32'hc19510c9, 32'hc1389160, 32'h42a39d39, 32'h424a702c, 32'h4218ad26, 32'hc2a86f3e};
test_label[195] = '{32'hc29b15fb};
test_output[195] = '{32'h431f599a};
/*############ DEBUG ############
test_input[1560:1567] = '{-77.5429338768, 8.71885454807, -18.6331957481, -11.5354917447, 81.8070786619, 50.6095422158, 38.169091451, -84.217269169};
test_label[195] = '{-77.5429338768};
test_output[195] = '{159.350012539};
############ END DEBUG ############*/
test_input[1568:1575] = '{32'hc1856d4e, 32'hc1cd1230, 32'hc2598b74, 32'hc2a16d6e, 32'h4271bd77, 32'h418c5a90, 32'hc2413e9b, 32'hc25d76b6};
test_label[196] = '{32'hc1856d4e};
test_output[196] = '{32'h429a3a0f};
/*############ DEBUG ############
test_input[1568:1575] = '{-16.6783716755, -25.6338812352, -54.3861842033, -80.713727059, 60.4350261564, 17.544219859, -48.3111381666, -55.3659273142};
test_label[196] = '{-16.6783716755};
test_output[196] = '{77.1133978319};
############ END DEBUG ############*/
test_input[1576:1583] = '{32'h4276c364, 32'h4290ab0e, 32'hc1667998, 32'hc1bcd526, 32'h42b963a2, 32'h42853aa2, 32'hc2b60380, 32'hc1fd68b5};
test_label[197] = '{32'hc1bcd526};
test_output[197] = '{32'h42e898eb};
/*############ DEBUG ############
test_input[1576:1583] = '{61.6908094685, 72.3340892915, -14.4046856197, -23.6040756468, 92.6945947849, 66.6145173618, -91.0068344787, -31.6761256799};
test_label[197] = '{-23.6040756468};
test_output[197] = '{116.298670433};
############ END DEBUG ############*/
test_input[1584:1591] = '{32'h4228b44a, 32'h4261047a, 32'h420e48ab, 32'hc284fb9b, 32'hc1e580c6, 32'hc1ab108c, 32'hc1f5624f, 32'h42c0aa75};
test_label[198] = '{32'h4228b44a};
test_output[198] = '{32'h4258a09f};
/*############ DEBUG ############
test_input[1584:1591] = '{42.1760653732, 56.2543711672, 35.5709663847, -66.4914164947, -28.6878785334, -21.3830800557, -30.6730016879, 96.3329224699};
test_label[198] = '{42.1760653732};
test_output[198] = '{54.1568570968};
############ END DEBUG ############*/
test_input[1592:1599] = '{32'hc213e393, 32'h41ccf33d, 32'h42843948, 32'h424432fc, 32'h424ba619, 32'hc1b1c63c, 32'hc2c1c299, 32'h42909179};
test_label[199] = '{32'h42909179};
test_output[199] = '{32'h3b0899df};
/*############ DEBUG ############
test_input[1592:1599] = '{-36.9722400915, 25.6187686101, 66.1118754455, 49.0497875527, 50.9122056572, -22.2217950291, -96.8800700698, 72.2841235801};
test_label[199] = '{72.2841235801};
test_output[199] = '{0.00208436670287};
############ END DEBUG ############*/
test_input[1600:1607] = '{32'h42a27dc7, 32'hc237fea6, 32'hc24591c4, 32'hc281d7af, 32'h42b171df, 32'hc2a5afb5, 32'h428f7e81, 32'h42006edf};
test_label[200] = '{32'hc237fea6};
test_output[200] = '{32'h4306b8be};
/*############ DEBUG ############
test_input[1600:1607] = '{81.2456593645, -45.9986803206, -49.3923475887, -64.9212569129, 88.7224065829, -82.8431761571, 71.7470805141, 32.1082717232};
test_label[200] = '{-45.9986803206};
test_output[200] = '{134.721652881};
############ END DEBUG ############*/
test_input[1608:1615] = '{32'h4228a9f6, 32'hc2c48594, 32'h42be7759, 32'h42b81471, 32'h409a80b9, 32'h42661ce9, 32'hc132f964, 32'hc2968342};
test_label[201] = '{32'h42b81471};
test_output[201] = '{32'h404eeff8};
/*############ DEBUG ############
test_input[1608:1615] = '{42.1659786834, -98.2608972835, 95.2331015789, 92.0399266584, 4.8282130138, 57.5282306753, -11.1858868503, -75.2563647353};
test_label[201] = '{92.0399266584};
test_output[201] = '{3.2333964412};
############ END DEBUG ############*/
test_input[1616:1623] = '{32'h4027c8c2, 32'hc214954c, 32'h41e9a858, 32'hc2b05b02, 32'h4295782f, 32'h42631980, 32'hc18abedf, 32'hc0871f22};
test_label[202] = '{32'hc0871f22};
test_output[202] = '{32'h429dea21};
/*############ DEBUG ############
test_input[1616:1623] = '{2.62162824984, -37.1457980533, 29.2071993689, -88.1777509184, 74.734736287, 56.7749018416, -17.3431981014, -4.22255050204};
test_label[202] = '{-4.22255050204};
test_output[202] = '{78.9572868049};
############ END DEBUG ############*/
test_input[1624:1631] = '{32'hc29f684c, 32'h42903dfe, 32'hc18efc5c, 32'hc2316973, 32'hc2c64256, 32'h41c2ddca, 32'hc2028939, 32'h4262f548};
test_label[203] = '{32'h41c2ddca};
test_output[203] = '{32'h423f0d17};
/*############ DEBUG ############
test_input[1624:1631] = '{-79.7037069169, 72.1210773285, -17.8732219949, -44.3529791221, -99.1295649776, 24.3582954032, -32.6340060736, 56.739531015};
test_label[203] = '{24.3582954032};
test_output[203] = '{47.7627821341};
############ END DEBUG ############*/
test_input[1632:1639] = '{32'h4025ab21, 32'h4262bf23, 32'hc2ab5298, 32'hc2b51428, 32'hc25ffb88, 32'h425e4707, 32'h41959020, 32'hc2ae74ad};
test_label[204] = '{32'h4262bf23};
test_output[204] = '{32'h3e90eb2b};
/*############ DEBUG ############
test_input[1632:1639] = '{2.58856982881, 56.6866569089, -85.6613142874, -90.5393645241, -55.9956359632, 55.5693625609, 18.6953728907, -87.2278804158};
test_label[204] = '{56.6866569089};
test_output[204] = '{0.283044176189};
############ END DEBUG ############*/
test_input[1640:1647] = '{32'hc2653f02, 32'h42ae6c03, 32'hc293736a, 32'hc24ae8a5, 32'h4242a6f7, 32'hc1791098, 32'h42af3ed1, 32'h42854925};
test_label[205] = '{32'hc293736a};
test_output[205] = '{32'h4321db3f};
/*############ DEBUG ############
test_input[1640:1647] = '{-57.3115319626, 87.2109635368, -73.7254209364, -50.7271925665, 48.6630508412, -15.5665511734, 87.6226907466, 66.6428612043};
test_label[205] = '{-73.7254209364};
test_output[205] = '{161.85643717};
############ END DEBUG ############*/
test_input[1648:1655] = '{32'h410e72e0, 32'hc1072aa5, 32'hc0f54f39, 32'hc2b1585f, 32'h423e497e, 32'h41cc88ca, 32'h42938cc7, 32'hc2810e02};
test_label[206] = '{32'h41cc88ca};
test_output[206] = '{32'h4240d529};
/*############ DEBUG ############
test_input[1648:1655] = '{8.90304530008, -8.4479111412, -7.66592073729, -88.6725971279, 47.5717687201, 25.5667923277, 73.7749546499, -64.5273590479};
test_label[206] = '{25.5667923277};
test_output[206] = '{48.2081623221};
############ END DEBUG ############*/
test_input[1656:1663] = '{32'hc27884c2, 32'h41925a8b, 32'hc27037da, 32'h429d128f, 32'hc29d1581, 32'hc28db08a, 32'hc24a8f7f, 32'hc29e9317};
test_label[207] = '{32'hc29d1581};
test_output[207] = '{32'h431d1408};
/*############ DEBUG ############
test_input[1656:1663] = '{-62.1296455973, 18.2942112728, -60.0545424921, 78.5362451729, -78.5419977246, -70.8448055426, -50.6401315896, -79.2872852632};
test_label[207] = '{-78.5419977246};
test_output[207] = '{157.078242898};
############ END DEBUG ############*/
test_input[1664:1671] = '{32'h424258cd, 32'hc251852d, 32'h423873ad, 32'hc049ef94, 32'hbf066e51, 32'h41ff08f1, 32'hc19d0e47, 32'hc1ef6896};
test_label[208] = '{32'hc251852d};
test_output[208] = '{32'h42ca1869};
/*############ DEBUG ############
test_input[1664:1671] = '{48.5867212355, -52.3800536726, 46.1129657562, -3.1552476424, -0.525120791554, 31.879365036, -19.6319715744, -29.9260678079};
test_label[208] = '{-52.3800536726};
test_output[208] = '{101.047679878};
############ END DEBUG ############*/
test_input[1672:1679] = '{32'h4229a43a, 32'hc2c36c38, 32'h42ad9d0d, 32'hc1b6aad0, 32'hc2c1f08f, 32'h3e3d8158, 32'h41c99815, 32'hc1b20470};
test_label[209] = '{32'h42ad9d0d};
test_output[209] = '{32'h80000000};
/*############ DEBUG ############
test_input[1672:1679] = '{42.4103764356, -97.7113648587, 86.8067425021, -22.8334042495, -96.969840035, 0.185063713066, 25.1992591451, -22.2521659804};
test_label[209] = '{86.8067425021};
test_output[209] = '{-0.0};
############ END DEBUG ############*/
test_input[1680:1687] = '{32'hc22e2160, 32'h4293777b, 32'h42a962e0, 32'h429b7705, 32'h428c9278, 32'hc1427213, 32'h4286127e, 32'hc2957847};
test_label[210] = '{32'h429b7705};
test_output[210] = '{32'h40dec58c};
/*############ DEBUG ############
test_input[1680:1687] = '{-43.5325944418, 73.7333589403, 84.6931124469, 77.7324636707, 70.2860721512, -12.15285024, 67.0361184381, -74.7349178417};
test_label[210] = '{77.7324636707};
test_output[210] = '{6.96161475306};
############ END DEBUG ############*/
test_input[1688:1695] = '{32'hc18010aa, 32'h425350be, 32'h41bcb0b4, 32'hc26aeab3, 32'h41e3951f, 32'hc2949dc5, 32'hc0d9ab72, 32'h420f3bd6};
test_label[211] = '{32'hc26aeab3};
test_output[211] = '{32'h42df1db8};
/*############ DEBUG ############
test_input[1688:1695] = '{-16.0081368408, 52.8288488004, 23.5862812095, -58.7291993401, 28.4478135793, -74.3081428695, -6.80217825329, 35.8084333273};
test_label[211] = '{-58.7291993401};
test_output[211] = '{111.558048181};
############ END DEBUG ############*/
test_input[1696:1703] = '{32'h42af0778, 32'hc29b938f, 32'h429342ef, 32'h428f08fe, 32'hc1efcabf, 32'h4292ddde, 32'hc29f28af, 32'h41d4c7d0};
test_label[212] = '{32'hc29b938f};
test_output[212] = '{32'h43254d84};
/*############ DEBUG ############
test_input[1696:1703] = '{87.5145910931, -77.788203329, 73.6307320355, 71.5175620902, -29.9739962658, 73.4333320049, -79.5794597081, 26.5975640722};
test_label[212] = '{-77.788203329};
test_output[212] = '{165.302796236};
############ END DEBUG ############*/
test_input[1704:1711] = '{32'h42768a19, 32'h4270a8ed, 32'h428dea11, 32'hc27fc596, 32'h42aa80d0, 32'hc292f332, 32'h4241b0a5, 32'h42750256};
test_label[213] = '{32'h428dea11};
test_output[213] = '{32'h4164b5fa};
/*############ DEBUG ############
test_input[1704:1711] = '{61.6348613583, 60.1649674615, 70.9571599552, -63.9429543306, 85.2515870277, -73.4749940169, 48.4225058863, 61.2522800285};
test_label[213] = '{70.9571599552};
test_output[213] = '{14.2944276921};
############ END DEBUG ############*/
test_input[1712:1719] = '{32'hc2948c54, 32'h42b7a5db, 32'h4208c335, 32'hc2c06876, 32'h42572426, 32'h426f3f2e, 32'hc25d603b, 32'h41e1db6e};
test_label[214] = '{32'h426f3f2e};
test_output[214] = '{32'h42000c89};
/*############ DEBUG ############
test_input[1712:1719] = '{-74.2740814592, 91.8239379932, 34.1906317328, -96.2040255887, 53.7853006063, 59.8116984226, -55.3439732616, 28.2321434505};
test_label[214] = '{59.8116984226};
test_output[214] = '{32.0122395706};
############ END DEBUG ############*/
test_input[1720:1727] = '{32'h4117b687, 32'hc1f4adff, 32'hc29825d0, 32'hc1c4f6b8, 32'h42ba11d3, 32'hc2a227ed, 32'h42ba52bc, 32'h42529275};
test_label[215] = '{32'h4117b687};
test_output[215] = '{32'h42a89f62};
/*############ DEBUG ############
test_input[1720:1727] = '{9.48206278753, -30.5849599534, -76.0738555937, -24.6204686601, 93.0348137756, -81.0779791434, 93.1615906535, 52.6430247435};
test_label[215] = '{9.48206278753};
test_output[215] = '{84.3112943107};
############ END DEBUG ############*/
test_input[1728:1735] = '{32'h423d862d, 32'h42a07dea, 32'h42b9ff70, 32'h4214ade9, 32'h41ade352, 32'hc26b9e8b, 32'hc2299d85, 32'h424cad88};
test_label[216] = '{32'hc2299d85};
test_output[216] = '{32'h43076719};
/*############ DEBUG ############
test_input[1728:1735] = '{47.381029684, 80.2459247762, 92.9989004434, 37.1698354891, 21.7359958303, -58.904825387, -42.4038284945, 51.1694651604};
test_label[216] = '{-42.4038284945};
test_output[216] = '{135.402731832};
############ END DEBUG ############*/
test_input[1736:1743] = '{32'h423a21e2, 32'hc22271fb, 32'h421ee24b, 32'hc28f9935, 32'hc2c212c9, 32'h40ad020d, 32'h428dde41, 32'h41ad1209};
test_label[217] = '{32'h40ad020d};
test_output[217] = '{32'h42830e20};
/*############ DEBUG ############
test_input[1736:1743] = '{46.5330905407, -40.6113092193, 39.7209883272, -71.7992315041, -97.0366863448, 5.4065004422, 70.934090173, 21.6338065505};
test_label[217] = '{5.4065004422};
test_output[217] = '{65.5275897308};
############ END DEBUG ############*/
test_input[1744:1751] = '{32'h40c48698, 32'h42ac40b6, 32'h42baf99f, 32'hc132547e, 32'hc2be6553, 32'h41ba8a8b, 32'hc1f1d366, 32'h42b2cc1b};
test_label[218] = '{32'h40c48698};
test_output[218] = '{32'h42aeba0a};
/*############ DEBUG ############
test_input[1744:1751] = '{6.14142981244, 86.1263847681, 93.4875439432, -11.1456281354, -95.1978970236, 23.3176475395, -30.2282215114, 89.3986422865};
test_label[218] = '{6.14142981244};
test_output[218] = '{87.3633576928};
############ END DEBUG ############*/
test_input[1752:1759] = '{32'h42611219, 32'h4283634a, 32'hc268a80e, 32'h402481f7, 32'h423caace, 32'h42348304, 32'hc2290e61, 32'hc238f087};
test_label[219] = '{32'h402481f7};
test_output[219] = '{32'h427c7e89};
/*############ DEBUG ############
test_input[1752:1759] = '{56.2676720914, 65.6939225615, -58.164115706, 2.57043241945, 47.1668012778, 45.127943354, -42.264043758, -46.2348886099};
test_label[219] = '{2.57043241945};
test_output[219] = '{63.1235707298};
############ END DEBUG ############*/
test_input[1760:1767] = '{32'hc188d42e, 32'hc22ae761, 32'h41625c90, 32'h4156f712, 32'hc2bb91cf, 32'h424628c0, 32'h42268020, 32'h42896466};
test_label[220] = '{32'hc22ae761};
test_output[220] = '{32'h42ded817};
/*############ DEBUG ############
test_input[1760:1767] = '{-17.1036031202, -42.7259564109, 14.1475985995, 13.4353203721, -93.7847814021, 49.539793347, 41.6251209642, 68.6960907772};
test_label[220] = '{-42.7259564109};
test_output[220] = '{111.422047193};
############ END DEBUG ############*/
test_input[1768:1775] = '{32'hc22f94c2, 32'h423b9306, 32'hc2025513, 32'hc177163e, 32'hc28f696c, 32'h42574278, 32'hc282dd5e, 32'hc1f472b2};
test_label[221] = '{32'hc1f472b2};
test_output[221] = '{32'h42a8be6a};
/*############ DEBUG ############
test_input[1768:1775] = '{-43.8952726034, 46.8935763233, -32.5830811218, -15.4429298752, -71.7058995251, 53.8149123169, -65.4323581776, -30.5560037309};
test_label[221] = '{-30.5560037309};
test_output[221] = '{84.3719020726};
############ END DEBUG ############*/
test_input[1776:1783] = '{32'h417579c7, 32'hc25d6c0c, 32'hc2c3aa7d, 32'h423c4e66, 32'h427a1c0e, 32'h418b5874, 32'hc0d56d1c, 32'h425bcb4a};
test_label[222] = '{32'hc2c3aa7d};
test_output[222] = '{32'h43205c63};
/*############ DEBUG ############
test_input[1776:1783] = '{15.3422308303, -55.3555148622, -97.8329827487, 47.076559509, 62.5273986401, 17.418189966, -6.66956919715, 54.9485237319};
test_label[222] = '{-97.8329827487};
test_output[222] = '{160.360892589};
############ END DEBUG ############*/
test_input[1784:1791] = '{32'h4266281a, 32'hc2aa17ac, 32'hc24d040d, 32'hc257f612, 32'hc2a92fcd, 32'hc193843a, 32'h414e4a36, 32'h423bede2};
test_label[223] = '{32'hc24d040d};
test_output[223] = '{32'h42d99617};
/*############ DEBUG ############
test_input[1784:1791] = '{57.5391625417, -85.0462327006, -51.2539554288, -53.9903022915, -84.5933638785, -18.4395628983, 12.8931177985, 46.9823058232};
test_label[223] = '{-51.2539554288};
test_output[223] = '{108.793143985};
############ END DEBUG ############*/
test_input[1792:1799] = '{32'hc29253fb, 32'h419fdb70, 32'h4167d7f2, 32'h42bdf463, 32'h42868981, 32'hc2b89af0, 32'hc21b82b0, 32'h42260d5e};
test_label[224] = '{32'h42260d5e};
test_output[224] = '{32'h4255db68};
/*############ DEBUG ############
test_input[1792:1799] = '{-73.1640278121, 19.9821480849, 14.4902210959, 94.977314623, 67.2685654771, -92.302609254, -38.8776257239, 41.5130525005};
test_label[224] = '{41.5130525005};
test_output[224] = '{53.4642621226};
############ END DEBUG ############*/
test_input[1800:1807] = '{32'h40afeb4b, 32'hc12cbfd2, 32'h42bd755e, 32'hc29b277c, 32'hc2c06a3f, 32'hc2a4ac01, 32'hc2940bae, 32'hc1f1673b};
test_label[225] = '{32'h42bd755e};
test_output[225] = '{32'h80000000};
/*############ DEBUG ############
test_input[1800:1807] = '{5.49747234977, -10.7968311608, 94.7292340028, -77.5771209131, -96.2075085189, -82.3359446973, -74.0228150666, -30.1754055763};
test_label[225] = '{94.7292340028};
test_output[225] = '{-0.0};
############ END DEBUG ############*/
test_input[1808:1815] = '{32'h42540123, 32'hc28d4290, 32'hc2918363, 32'hc116d966, 32'hc21bdb5c, 32'h42255581, 32'h42767dc6, 32'h42310f3c};
test_label[226] = '{32'h42767dc6};
test_output[226] = '{32'h393ceac5};
/*############ DEBUG ############
test_input[1808:1815] = '{53.0011112405, -70.6300012085, -72.7566161247, -9.42807616889, -38.9642166583, 41.3334987843, 61.6228258217, 44.2648773325};
test_label[226] = '{61.6228258217};
test_output[226] = '{0.000180165361296};
############ END DEBUG ############*/
test_input[1816:1823] = '{32'h421bee73, 32'h428b51c5, 32'h4286bb33, 32'hc29e3c80, 32'h41071567, 32'hc2bbb288, 32'hc13ed154, 32'hc2bae10e};
test_label[227] = '{32'hc2bae10e};
test_output[227] = '{32'h43233203};
/*############ DEBUG ############
test_input[1816:1823] = '{38.9828606458, 69.6597080111, 67.3656222851, -79.1181629792, 8.44272541871, -93.8486912902, -11.9261050486, -93.4395622365};
test_label[227] = '{-93.4395622365};
test_output[227] = '{163.195356089};
############ END DEBUG ############*/
test_input[1824:1831] = '{32'hc2b38f71, 32'h42b5bd9c, 32'h41d87eff, 32'hc1f0d24a, 32'h41cb22f4, 32'h3d6fccd7, 32'h42b3b106, 32'h417f761a};
test_label[228] = '{32'h41d87eff};
test_output[228] = '{32'h42803ae6};
/*############ DEBUG ############
test_input[1824:1831] = '{-89.7801587648, 90.8703343715, 27.062009574, -30.1026810603, 25.3920665276, 0.0585449581243, 89.845746558, 15.9663332795};
test_label[228] = '{27.062009574};
test_output[228] = '{64.1150330098};
############ END DEBUG ############*/
test_input[1832:1839] = '{32'h41163268, 32'hc239a79a, 32'h423fe1ba, 32'h422cd4ce, 32'h424a5f10, 32'h42884347, 32'h409aa767, 32'hc185986c};
test_label[229] = '{32'h422cd4ce};
test_output[229] = '{32'h41c7637e};
/*############ DEBUG ############
test_input[1832:1839] = '{9.38730594036, -46.4136723489, 47.9704371528, 43.2078164407, 50.5928329869, 68.1313975151, 4.83293491686, -16.6994255352};
test_label[229] = '{43.2078164407};
test_output[229] = '{24.9235811003};
############ END DEBUG ############*/
test_input[1840:1847] = '{32'h42881a13, 32'hc2343bfd, 32'hc298bfd6, 32'h42962d71, 32'hc2991d2d, 32'hc194af16, 32'h42aeb44c, 32'hc247f864};
test_label[230] = '{32'hc194af16};
test_output[230] = '{32'h42d3e012};
/*############ DEBUG ############
test_input[1840:1847] = '{68.0509249441, -45.0585839394, -76.3746772271, 75.0887514976, -76.5569864758, -18.5854920835, 87.3521392793, -49.9925687767};
test_label[230] = '{-18.5854920835};
test_output[230] = '{105.937636088};
############ END DEBUG ############*/
test_input[1848:1855] = '{32'hc1f6a1cb, 32'h428ef469, 32'h428ecf38, 32'hc2bc3822, 32'h41bb62bb, 32'h42a0d2c4, 32'h42350f6c, 32'hc2c2001d};
test_label[231] = '{32'h428ef469};
test_output[231] = '{32'h410ef3e4};
/*############ DEBUG ############
test_input[1848:1855] = '{-30.8290001969, 71.4773631413, 71.4047222286, -94.1096307625, 23.4232080237, 80.4116528707, 45.2650585178, -97.0002236517};
test_label[231] = '{71.4773631413};
test_output[231] = '{8.93454404606};
############ END DEBUG ############*/
test_input[1856:1863] = '{32'hc262d8f8, 32'h426c17c8, 32'h42b62971, 32'hc16e46b2, 32'hc1ada43a, 32'hc1a36344, 32'h428ef499, 32'hc2a035bd};
test_label[232] = '{32'hc16e46b2};
test_output[232] = '{32'h42d3f247};
/*############ DEBUG ############
test_input[1856:1863] = '{-56.7118819804, 59.0232242023, 91.0809364816, -14.8922599829, -21.7051879467, -20.4234690952, 71.4777260665, -80.1049602223};
test_label[232] = '{-14.8922599829};
test_output[232] = '{105.973196468};
############ END DEBUG ############*/
test_input[1864:1871] = '{32'hc2a04554, 32'h422bcffb, 32'h424dea54, 32'hc0bea9ec, 32'hc25eff0c, 32'h424492ea, 32'h41bb0fe4, 32'h42a2bf4f};
test_label[233] = '{32'h41bb0fe4};
test_output[233] = '{32'h4267f6ad};
/*############ DEBUG ############
test_input[1864:1871] = '{-80.1354031345, 42.9531052156, 51.4788350327, -5.95824228625, -55.7490683158, 49.1434705689, 23.3827588724, 81.3736513615};
test_label[233] = '{23.3827588724};
test_output[233] = '{57.9908924892};
############ END DEBUG ############*/
test_input[1872:1879] = '{32'h4286d211, 32'h41c778cd, 32'h41aa89c0, 32'h42a4eb80, 32'hc2a75886, 32'hc01d8126, 32'hc1bf6d56, 32'h426213c7};
test_label[234] = '{32'h42a4eb80};
test_output[234] = '{32'h349c4657};
/*############ DEBUG ############
test_input[1872:1879] = '{67.4102877833, 24.9339840999, 21.3172613916, 82.4599586792, -83.6728938179, -2.46100763803, -23.928386474, 56.5193122364};
test_label[234] = '{82.4599586792};
test_output[234] = '{2.91084446945e-07};
############ END DEBUG ############*/
test_input[1880:1887] = '{32'hc10a3ed0, 32'hc164cd5c, 32'hc23f9c57, 32'h40b3e5a1, 32'hc2b75eb5, 32'h41967cb5, 32'h4295379a, 32'h42c386e0};
test_label[235] = '{32'h4295379a};
test_output[235] = '{32'h41b93d1a};
/*############ DEBUG ############
test_input[1880:1887] = '{-8.64033475268, -14.3001366838, -47.9026743361, 5.62178089623, -91.6849761735, 18.8108914729, 74.6085933156, 97.763427846};
test_label[235] = '{74.6085933156};
test_output[235] = '{23.1548345305};
############ END DEBUG ############*/
test_input[1888:1895] = '{32'hc299ebb9, 32'h42b4d134, 32'hc197a0ee, 32'hc093b006, 32'h42ae52ae, 32'h4226da8d, 32'h428fff85, 32'hc2bcb68d};
test_label[236] = '{32'h42b4d134};
test_output[236] = '{32'h3d1c4260};
/*############ DEBUG ############
test_input[1888:1895] = '{-76.9603940989, 90.4085981701, -18.9535798421, -4.61523736471, 87.1614836162, 41.7134301047, 71.9990606233, -94.3565420392};
test_label[236] = '{90.4085981701};
test_output[236] = '{0.0381492358665};
############ END DEBUG ############*/
test_input[1896:1903] = '{32'h4287e47a, 32'hbff7cd1e, 32'hc24d8b03, 32'hc1e406a1, 32'h429238c9, 32'hc19317b6, 32'hc148e4f4, 32'hc2ada9dc};
test_label[237] = '{32'h429238c9};
test_output[237] = '{32'h3bbabc25};
/*############ DEBUG ############
test_input[1896:1903] = '{67.9462433744, -1.93594718873, -51.3857527817, -28.503236979, 73.11091022, -18.3865768467, -12.5558969404, -86.8317580005};
test_label[237] = '{73.11091022};
test_output[237] = '{0.00569869802023};
############ END DEBUG ############*/
test_input[1904:1911] = '{32'h416eda61, 32'h42c29f0a, 32'hc09c1e25, 32'h42213072, 32'h42b05b53, 32'h41e8d381, 32'hc2a5ddbc, 32'h42867fa7};
test_label[238] = '{32'h416eda61};
test_output[238] = '{32'h42a4c3cc};
/*############ DEBUG ############
test_input[1904:1911] = '{14.9283149924, 97.3106196353, -4.87867990333, 40.2973090619, 88.1783650697, 29.1032726713, -82.9330749684, 67.2493177947};
test_label[238] = '{14.9283149924};
test_output[238] = '{82.3824127586};
############ END DEBUG ############*/
test_input[1912:1919] = '{32'h3fb1b83d, 32'hc2152285, 32'hc18d98eb, 32'h4284f17c, 32'h400ad7ef, 32'hc2081345, 32'h4287eb55, 32'h429a0452};
test_label[239] = '{32'h4284f17c};
test_output[239] = '{32'h41289743};
/*############ DEBUG ############
test_input[1912:1919] = '{1.38843500196, -37.2837111154, -17.6996662252, 66.4716509105, 2.16942944663, -34.018818696, 67.9596308605, 77.00843564};
test_label[239] = '{66.4716509105};
test_output[239] = '{10.5369287925};
############ END DEBUG ############*/
test_input[1920:1927] = '{32'hc0d6a054, 32'h42b14432, 32'hc19a80ee, 32'h42a4f768, 32'hc2729ca0, 32'h40fc5ff5, 32'h42784b36, 32'h4185a729};
test_label[240] = '{32'hc2729ca0};
test_output[240] = '{32'h431549cc};
/*############ DEBUG ############
test_input[1920:1927] = '{-6.70707111167, 88.6331914239, -19.3129532313, 82.4832149291, -60.6529536407, 7.88671336476, 62.0734469961, 16.7066215436};
test_label[240] = '{-60.6529536407};
test_output[240] = '{149.288276324};
############ END DEBUG ############*/
test_input[1928:1935] = '{32'h42af7ca6, 32'hc21b0e5f, 32'h4263711d, 32'hc2ab99f8, 32'h425909a8, 32'hc23f546f, 32'hc1cbb5bd, 32'hc2a2a35d};
test_label[241] = '{32'hc2a2a35d};
test_output[241] = '{32'h43291002};
/*############ DEBUG ############
test_input[1928:1935] = '{87.7434554884, -38.7640324984, 56.8604633323, -85.8007187905, 54.2594310039, -47.8324550196, -25.4637395804, -81.319071522};
test_label[241] = '{-81.319071522};
test_output[241] = '{169.06252701};
############ END DEBUG ############*/
test_input[1936:1943] = '{32'h41e5c630, 32'hc1aee548, 32'h41c316e5, 32'h4268d283, 32'hc185e15e, 32'h426fbc2d, 32'h40cd157a, 32'hc2805f96};
test_label[242] = '{32'h41e5c630};
test_output[242] = '{32'h41fb00fa};
/*############ DEBUG ############
test_input[1936:1943] = '{28.7217719387, -21.8619535986, 24.386178849, 58.2055770184, -16.7350419451, 59.933765535, 6.40887170303, -64.1866947601};
test_label[242] = '{28.7217719387};
test_output[242] = '{31.375477032};
############ END DEBUG ############*/
test_input[1944:1951] = '{32'h42c12c02, 32'h42830349, 32'hc20af60f, 32'h41a2f344, 32'h423c1b62, 32'h3f1f57d4, 32'hc2861d11, 32'h428b574d};
test_label[243] = '{32'h428b574d};
test_output[243] = '{32'h41d752d6};
/*############ DEBUG ############
test_input[1944:1951] = '{96.5859538759, 65.506419157, -34.7402901744, 20.3687825362, 47.0267397979, 0.622433893826, -67.0567690503, 69.6705069269};
test_label[243] = '{69.6705069269};
test_output[243] = '{26.915446949};
############ END DEBUG ############*/
test_input[1952:1959] = '{32'h419699e7, 32'h42c1ad53, 32'h413bfe37, 32'hc2afa41b, 32'h423bd3f9, 32'h423f99e9, 32'hc2869a6c, 32'hc2956088};
test_label[244] = '{32'hc2869a6c};
test_output[244] = '{32'h432423e0};
/*############ DEBUG ############
test_input[1952:1959] = '{18.8251471308, 96.8385267848, 11.749564642, -87.8205207737, 46.9570055756, 47.9003010558, -67.3016047048, -74.688537326};
test_label[244] = '{-67.3016047048};
test_output[244] = '{164.14013149};
############ END DEBUG ############*/
test_input[1960:1967] = '{32'h41d81cd8, 32'hc2b7556d, 32'hc0f6572a, 32'hc28d2b98, 32'hc2881d94, 32'hc278abc1, 32'h4216529d, 32'h41fbbfbf};
test_label[245] = '{32'hc28d2b98};
test_output[245] = '{32'h42d8560c};
/*############ DEBUG ############
test_input[1960:1967] = '{27.0140843879, -91.6668485986, -7.69814034923, -70.5851453958, -68.057767185, -62.1677272138, 37.5806768276, 31.468626917};
test_label[245] = '{-70.5851453958};
test_output[245] = '{108.16806148};
############ END DEBUG ############*/
test_input[1968:1975] = '{32'hc27e3f16, 32'hc2071a56, 32'hc28b5773, 32'hc296c31e, 32'h41b88d56, 32'hc267a0ee, 32'h41a764a8, 32'h4203fc34};
test_label[246] = '{32'h4203fc34};
test_output[246] = '{32'h3864c15c};
/*############ DEBUG ############
test_input[1968:1975] = '{-63.5616064723, -33.7757182663, -69.6708024589, -75.3810901129, 23.0690114427, -57.9071561908, 20.924148525, 32.9962910134};
test_label[246] = '{32.9962910134};
test_output[246] = '{5.45395165477e-05};
############ END DEBUG ############*/
test_input[1976:1983] = '{32'hc240e299, 32'h4282fac6, 32'hc1d1f408, 32'h426a1afb, 32'hc2a27968, 32'h428c864d, 32'h414e04a9, 32'h3d73ad29};
test_label[247] = '{32'hc240e299};
test_output[247] = '{32'h42ecfbeb};
/*############ DEBUG ############
test_input[1976:1983] = '{-48.2212876253, 65.4897910305, -26.2441555595, 58.5263494364, -81.2371242402, 70.2623058491, 12.8761372812, 0.0594913097799};
test_label[247] = '{-48.2212876253};
test_output[247] = '{118.492024911};
############ END DEBUG ############*/
test_input[1984:1991] = '{32'hc1e089bd, 32'hc294cf7b, 32'h426be6b8, 32'h428ef850, 32'h429655a7, 32'h41f57772, 32'h411cdb8f, 32'h42372a46};
test_label[248] = '{32'h411cdb8f};
test_output[248] = '{32'h4282c6ef};
/*############ DEBUG ############
test_input[1984:1991] = '{-28.0672551107, -74.4052352342, 58.9753099643, 71.484984641, 75.1672898451, 30.6833234363, 9.80360364663, 45.7912826455};
test_label[248] = '{9.80360364663};
test_output[248] = '{65.3885397646};
############ END DEBUG ############*/
test_input[1992:1999] = '{32'h423ddc22, 32'hc213847d, 32'h42bab79e, 32'h424c4aef, 32'h41329cf0, 32'h4184ba68, 32'h4218a774, 32'hc2b4c215};
test_label[249] = '{32'h42bab79e};
test_output[249] = '{32'h80000000};
/*############ DEBUG ############
test_input[1992:1999] = '{47.4649751784, -36.8793840773, 93.3586275213, 51.0731777543, 11.1633147613, 16.5910185075, 38.1635269317, -90.3790636646};
test_label[249] = '{93.3586275213};
test_output[249] = '{-0.0};
############ END DEBUG ############*/
test_input[2000:2007] = '{32'h4246c688, 32'h428ddefb, 32'h41bc7325, 32'h42be5281, 32'hc2b7b25e, 32'h42a938bd, 32'h425180c8, 32'hc1487087};
test_label[250] = '{32'hc1487087};
test_output[250] = '{32'h42d76095};
/*############ DEBUG ############
test_input[2000:2007] = '{49.6938796672, 70.9355070339, 23.5562231075, 95.1611387436, -91.8483751076, 84.6108146986, 52.3757610862, -12.5274726968};
test_label[250] = '{-12.5274726968};
test_output[250] = '{107.688637625};
############ END DEBUG ############*/
test_input[2008:2015] = '{32'hc2a3a91f, 32'hc2548ddf, 32'h42b13d4f, 32'hc2be5c36, 32'hc2360e88, 32'hc27beb0e, 32'h41a8f354, 32'h4180cc1d};
test_label[251] = '{32'hc27beb0e};
test_output[251] = '{32'h4317996b};
/*############ DEBUG ############
test_input[2008:2015] = '{-81.8303161729, -53.1385470224, 88.6197419845, -95.1801016759, -45.5141893165, -62.9795441193, 21.1188122176, 16.0996639895};
test_label[251] = '{-62.9795441193};
test_output[251] = '{151.599286104};
############ END DEBUG ############*/
test_input[2016:2023] = '{32'hc22345e7, 32'hc2583249, 32'hc2995911, 32'hc1817303, 32'hc282fb46, 32'h4258dab9, 32'hc20586cc, 32'h41d49f47};
test_label[252] = '{32'hc1817303};
test_output[252] = '{32'h428cca1d};
/*############ DEBUG ############
test_input[2016:2023] = '{-40.8182637288, -54.0491084069, -76.673957993, -16.1811583064, -65.4907654899, 54.2135963906, -33.3816381398, 26.5777725871};
test_label[252] = '{-16.1811583064};
test_output[252] = '{70.394754697};
############ END DEBUG ############*/
test_input[2024:2031] = '{32'hc2b0b9e3, 32'hc2c3ffeb, 32'h42187318, 32'h42310ff4, 32'h412eb972, 32'hc1d06246, 32'h4212df7c, 32'hc2925be5};
test_label[253] = '{32'hc1d06246};
test_output[253] = '{32'h428ca1e7};
/*############ DEBUG ############
test_input[2024:2031] = '{-88.3630589963, -97.9998377195, 38.1123970823, 44.2655808745, 10.9202745996, -26.0479849098, 36.7182468346, -73.1794831783};
test_label[253] = '{-26.0479849098};
test_output[253] = '{70.3162164828};
############ END DEBUG ############*/
test_input[2032:2039] = '{32'h41a40f22, 32'h4223a33f, 32'hc249c168, 32'h40bb817f, 32'h4215ae14, 32'hc217f2e9, 32'hc296c792, 32'h421208fc};
test_label[254] = '{32'h4215ae14};
test_output[254] = '{32'h40620124};
/*############ DEBUG ############
test_input[2032:2039] = '{20.5073881177, 40.9094207589, -50.4388736398, 5.85955758081, 37.4199990173, -37.9872153923, -75.3897866298, 36.5087738355};
test_label[254] = '{37.4199990173};
test_output[254] = '{3.5313195566};
############ END DEBUG ############*/
test_input[2040:2047] = '{32'h42ac7d68, 32'hc28ed75d, 32'h414d302c, 32'h42912594, 32'hc191949c, 32'hc1a3684c, 32'h41a40fbe, 32'h41d919a2};
test_label[255] = '{32'h41d919a2};
test_output[255] = '{32'h426c6dff};
/*############ DEBUG ############
test_input[2040:2047] = '{86.2449356206, -71.4206351246, 12.8242605519, 72.5733944617, -18.1975622716, -20.4259259083, 20.5076857647, 27.1375169644};
test_label[255] = '{27.1375169644};
test_output[255] = '{59.1074198111};
############ END DEBUG ############*/
test_input[2048:2055] = '{32'hc144eee3, 32'h4294fe0a, 32'hc139a1c0, 32'h42c45275, 32'h41c0d08a, 32'hc2149e44, 32'hc1f97ff4, 32'hc203d419};
test_label[256] = '{32'hc139a1c0};
test_output[256] = '{32'h42db86ad};
/*############ DEBUG ############
test_input[2048:2055] = '{-12.3083215403, 74.496166725, -11.6019893105, 98.1610504993, 24.1018248622, -37.1545565708, -31.1874768751, -32.9571276961};
test_label[256] = '{-11.6019893105};
test_output[256] = '{109.76303981};
############ END DEBUG ############*/
test_input[2056:2063] = '{32'hc225da39, 32'hc2ace7c2, 32'hc200419c, 32'h422f1648, 32'hc28c9871, 32'hc226d7b4, 32'h4287bcd8, 32'h4197e2f1};
test_label[257] = '{32'h422f1648};
test_output[257] = '{32'h41c0c6d1};
/*############ DEBUG ############
test_input[2056:2063] = '{-41.4631067619, -86.452652906, -32.0640733502, 43.7717577971, -70.2977384114, -41.7106464808, 67.8688352623, 18.985810664};
test_label[257] = '{43.7717577971};
test_output[257] = '{24.0970774652};
############ END DEBUG ############*/
test_input[2064:2071] = '{32'hc1dd615f, 32'hc212ed8f, 32'hc2ae6c46, 32'hc152ad1b, 32'hc2c375c7, 32'hc2c5a1f2, 32'hbe95d7c6, 32'hc11c71ad};
test_label[258] = '{32'hbe95d7c6};
test_output[258] = '{32'h38a4b35b};
/*############ DEBUG ############
test_input[2064:2071] = '{-27.6725453855, -36.7319918321, -87.2114682914, -13.1672624441, -97.7300345914, -98.8163021224, -0.292661850916, -9.77775306443};
test_label[258] = '{-0.292661850916};
test_output[258] = '{7.85353693372e-05};
############ END DEBUG ############*/
test_input[2072:2079] = '{32'h4293fbe0, 32'hc2c58e3a, 32'hc1c7a2ef, 32'h42307612, 32'h42aa97f5, 32'hc292e9ff, 32'hc281613f, 32'h40b46f44};
test_label[259] = '{32'h4293fbe0};
test_output[259] = '{32'h4134e0b5};
/*############ DEBUG ############
test_input[2072:2079] = '{73.9919400425, -98.7777872214, -24.9545575086, 44.1153031365, 85.296787778, -73.4570245409, -64.6899343329, 5.63858235845};
test_label[259] = '{73.9919400425};
test_output[259] = '{11.3048600485};
############ END DEBUG ############*/
test_input[2080:2087] = '{32'hc20362c6, 32'hc2918e17, 32'h4275cfd2, 32'h4275f331, 32'h424106e9, 32'h409d1985, 32'hc214f590, 32'h4236812c};
test_label[260] = '{32'hc20362c6};
test_output[260] = '{32'h42be051c};
/*############ DEBUG ############
test_input[2080:2087] = '{-32.8464602468, -72.7775203443, 61.4529494519, 61.4874903327, 48.2567483914, 4.90936498667, -37.2398057942, 45.6261435682};
test_label[260] = '{-32.8464602468};
test_output[260] = '{95.0099774248};
############ END DEBUG ############*/
test_input[2088:2095] = '{32'hc1cd3088, 32'h41fa6919, 32'h4240cad0, 32'hbf93a47f, 32'h41a35017, 32'h41a55a92, 32'hc23de04e, 32'hc18b6cbe};
test_label[261] = '{32'h41a55a92};
test_output[261] = '{32'h41dc3b0f};
/*############ DEBUG ############
test_input[2088:2095] = '{-25.6486976825, 31.3013164331, 48.1980604071, -1.1534575375, 20.4141068194, 20.6692240424, -47.4690471355, -17.428097303};
test_label[261] = '{20.6692240424};
test_output[261] = '{27.5288364106};
############ END DEBUG ############*/
test_input[2096:2103] = '{32'h426e808c, 32'hc27aa7a5, 32'h4298114e, 32'hc2c3dd50, 32'hc20c5e35, 32'hc20e4125, 32'hc29f42d4, 32'hc267f984};
test_label[262] = '{32'hc27aa7a5};
test_output[262] = '{32'h430ab290};
/*############ DEBUG ############
test_input[2096:2103] = '{59.6255334121, -62.6637145979, 76.0337993709, -97.9322483692, -35.0919987451, -35.563618379, -79.6305224434, -57.9936690284};
test_label[262] = '{-62.6637145979};
test_output[262] = '{138.697514044};
############ END DEBUG ############*/
test_input[2104:2111] = '{32'h41218646, 32'hc17f7d9b, 32'hc19a0349, 32'h419aa8b9, 32'h41cdb744, 32'h421683fb, 32'hc2bc6da2, 32'hc2096057};
test_label[263] = '{32'h421683fb};
test_output[263] = '{32'h36e0f815};
/*############ DEBUG ############
test_input[2104:2111] = '{10.0952816762, -15.9681653855, -19.2516042393, 19.3323840155, 25.7144848342, 37.6288883526, -94.2141253555, -34.3440835977};
test_label[263] = '{37.6288883526};
test_output[263] = '{6.70460087314e-06};
############ END DEBUG ############*/
test_input[2112:2119] = '{32'hc29e4c0d, 32'h420027f6, 32'h41bd3a4d, 32'h42a9e632, 32'h4279bbe9, 32'hc18ed357, 32'hc2839d85, 32'h4229f5e9};
test_label[264] = '{32'h41bd3a4d};
test_output[264] = '{32'h42752f3d};
/*############ DEBUG ############
test_input[2112:2119] = '{-79.1485387975, 32.0390228196, 23.6534676439, 84.949598588, 62.4335070465, -17.8531934969, -65.807658205, 42.4901461912};
test_label[264] = '{23.6534676439};
test_output[264] = '{61.2961309444};
############ END DEBUG ############*/
test_input[2120:2127] = '{32'hc2669066, 32'hc28b002d, 32'h4251e289, 32'h4231975d, 32'hc2bd4b0d, 32'h424f0eb3, 32'hc24ee183, 32'hc20cc82e};
test_label[265] = '{32'h4251e289};
test_output[265] = '{32'h3ecd5fa1};
/*############ DEBUG ############
test_input[2120:2127] = '{-57.6410145772, -69.5003411304, 52.4712262494, 44.3978173542, -94.6465828627, 51.7643554749, -51.7202270598, -35.1954896727};
test_label[265] = '{52.4712262494};
test_output[265] = '{0.401120210331};
############ END DEBUG ############*/
test_input[2128:2135] = '{32'hc112872e, 32'hc083b485, 32'hc277df86, 32'h404d3b20, 32'h4282d328, 32'h427161c8, 32'h41c26860, 32'h4136fd4f};
test_label[266] = '{32'h4282d328};
test_output[266] = '{32'h3bcdd910};
/*############ DEBUG ############
test_input[2128:2135] = '{-9.15800253663, -4.1157861441, -61.9682858834, 3.2067337441, 65.4124153434, 60.3454877907, 24.3009634264, 11.4368430797};
test_label[266] = '{65.4124153434};
test_output[266] = '{0.00628197921424};
############ END DEBUG ############*/
test_input[2136:2143] = '{32'h41a0af8e, 32'hc214903b, 32'h424df63c, 32'h428bae76, 32'h42a0513e, 32'h4201bef5, 32'hc28c432c, 32'h42197c71};
test_label[267] = '{32'hc28c432c};
test_output[267] = '{32'h43164a37};
/*############ DEBUG ############
test_input[2136:2143] = '{20.0857199531, -37.1408490305, 51.4904640794, 69.8407443355, 80.1586775792, 32.4364828482, -70.1311980873, 38.3715260304};
test_label[267] = '{-70.1311980873};
test_output[267] = '{150.289908701};
############ END DEBUG ############*/
test_input[2144:2151] = '{32'hc23f76aa, 32'hc2a95cb6, 32'hc28ef5a8, 32'h410d3b89, 32'h42958f28, 32'h428f7c31, 32'h42483171, 32'hc291b519};
test_label[268] = '{32'hc28ef5a8};
test_output[268] = '{32'h43124e67};
/*############ DEBUG ############
test_input[2144:2151] = '{-47.8658818877, -84.6810764574, -71.4798001365, 8.82703483294, 74.7795984647, 71.7425607099, 50.0482831723, -72.8537052071};
test_label[268] = '{-71.4798001365};
test_output[268] = '{146.306260048};
############ END DEBUG ############*/
test_input[2152:2159] = '{32'hc2c51a97, 32'h42b98ce5, 32'h42c4f73b, 32'hc276d6f4, 32'h41e4ae1f, 32'hc284544d, 32'hc2955992, 32'h41083aad};
test_label[269] = '{32'h42b98ce5};
test_output[269] = '{32'h40b6c089};
/*############ DEBUG ############
test_input[2152:2159] = '{-98.5519313516, 92.7751853445, 98.4828732368, -61.709916558, 28.5850208773, -66.164647821, -74.6749398141, 8.51432475982};
test_label[269] = '{92.7751853445};
test_output[269] = '{5.71100273272};
############ END DEBUG ############*/
test_input[2160:2167] = '{32'h42737ed1, 32'h423bc7e0, 32'hc030bde3, 32'h412e703e, 32'h40c47161, 32'h4190429f, 32'h42bf0536, 32'hc21fc90a};
test_label[270] = '{32'h42bf0536};
test_output[270] = '{32'h26800000};
/*############ DEBUG ############
test_input[2160:2167] = '{60.8738455018, 46.9451919806, -2.76158973481, 10.902402859, 6.13884009561, 18.0325306869, 95.510178562, -39.9463255171};
test_label[270] = '{95.510178562};
test_output[270] = '{8.881784197e-16};
############ END DEBUG ############*/
test_input[2168:2175] = '{32'h3eb38c9e, 32'hc013b32e, 32'h419d84b6, 32'h42a78b12, 32'h41fb3fa7, 32'hc287e05b, 32'hc2302219, 32'h42c00221};
test_label[271] = '{32'h41fb3fa7};
test_output[271] = '{32'h42813238};
/*############ DEBUG ############
test_input[2168:2175] = '{0.350682209079, -2.30781131829, 19.6898008536, 83.7716203961, 31.4060808537, -67.9381971898, -44.0332987997, 96.0041562771};
test_label[271] = '{31.4060808537};
test_output[271] = '{64.5980802928};
############ END DEBUG ############*/
test_input[2176:2183] = '{32'h42ab3ef0, 32'h42b02138, 32'h42985001, 32'h427b906d, 32'h42b5e7f2, 32'h427eb508, 32'h410a55b1, 32'h4267222b};
test_label[272] = '{32'h42b02138};
test_output[272] = '{32'h403c9a06};
/*############ DEBUG ############
test_input[2176:2183] = '{85.6229214392, 88.0648769377, 76.1562562068, 62.8910393372, 90.9530148729, 63.6767879537, 8.6459208, 57.783365832};
test_label[272] = '{88.0648769377};
test_output[272] = '{2.94690086065};
############ END DEBUG ############*/
test_input[2184:2191] = '{32'hc21127a2, 32'h42076ec5, 32'hc13e2999, 32'h425cc68a, 32'hc29b4c22, 32'hc2615eac, 32'h41e4e164, 32'hc13ae708};
test_label[273] = '{32'hc13ae708};
test_output[273] = '{32'h4285c026};
/*############ DEBUG ############
test_input[2184:2191] = '{-36.2887026279, 33.8581723432, -11.8851557597, 55.1938875201, -77.6486944655, -56.3424515909, 28.6100547628, -11.6814039228};
test_label[273] = '{-11.6814039228};
test_output[273] = '{66.8752914434};
############ END DEBUG ############*/
test_input[2192:2199] = '{32'hc2bbcfcd, 32'hc001aeb9, 32'h4233bfc2, 32'hc2aa4463, 32'h42a4e419, 32'h3f705e44, 32'hc27317b3, 32'hc255319b};
test_label[274] = '{32'hc2aa4463};
test_output[274] = '{32'h4327943e};
/*############ DEBUG ############
test_input[2192:2199] = '{-93.9058647004, -2.02628925053, 44.9372622691, -85.1335679728, 82.4455064399, 0.938938383792, -60.7731429201, -53.2984442126};
test_label[274] = '{-85.1335679728};
test_output[274] = '{167.579074413};
############ END DEBUG ############*/
test_input[2200:2207] = '{32'h427a5cfd, 32'hc2a38a89, 32'h42803301, 32'h42166cc8, 32'hc1f00721, 32'h429dd06b, 32'hc21e7814, 32'h4209b600};
test_label[275] = '{32'hc1f00721};
test_output[275] = '{32'h42d9d234};
/*############ DEBUG ############
test_input[2200:2207] = '{62.5908100137, -81.7705735347, 64.0996202714, 37.6062303817, -30.0034810832, 78.9070691798, -39.617264681, 34.4277339084};
test_label[275] = '{-30.0034810832};
test_output[275] = '{108.910550716};
############ END DEBUG ############*/
test_input[2208:2215] = '{32'h4291f749, 32'hc2b5c3cd, 32'hc2339fbe, 32'h4190d4aa, 32'h40309192, 32'hc2c6234c, 32'h423b7355, 32'hc2585980};
test_label[276] = '{32'h4291f749};
test_output[276] = '{32'h2c9f6100};
/*############ DEBUG ############
test_input[2208:2215] = '{72.9829796454, -90.8824255774, -44.9059998438, 18.1038395073, 2.75888479112, -99.0689416119, 46.8626293196, -54.0874022575};
test_label[276] = '{72.9829796454};
test_output[276] = '{4.52982096278e-12};
############ END DEBUG ############*/
test_input[2216:2223] = '{32'hc24cc87c, 32'h423ae2ba, 32'hc23e8e21, 32'h42a38378, 32'hc1fe8b64, 32'h416313f3, 32'h40408cbb, 32'hc2c58f6a};
test_label[277] = '{32'hc24cc87c};
test_output[277] = '{32'h4304f3db};
/*############ DEBUG ############
test_input[2216:2223] = '{-51.1957853086, 46.7214130005, -47.6387982781, 81.756776072, -31.818061921, 14.1923702529, 3.00858961663, -98.780109332};
test_label[277] = '{-51.1957853086};
test_output[277] = '{132.952561381};
############ END DEBUG ############*/
test_input[2224:2231] = '{32'h419b6462, 32'hc28ad1c3, 32'h424e8872, 32'h41963cc4, 32'hc1659c47, 32'hc29e3cce, 32'hc298b374, 32'hc134a1ab};
test_label[278] = '{32'h419b6462};
test_output[278] = '{32'h4200d641};
/*############ DEBUG ############
test_input[2224:2231] = '{19.4240151004, -69.4096932221, 51.6332461396, 18.7796712891, -14.3506540725, -79.1187605772, -76.3504928621, -11.2894693275};
test_label[278] = '{19.4240151004};
test_output[278] = '{32.2092310392};
############ END DEBUG ############*/
test_input[2232:2239] = '{32'h4117e3b7, 32'hc2c48be1, 32'hc2a2e484, 32'h4299f737, 32'hc255777e, 32'hc262d097, 32'hc2b2293c, 32'h42a87cf8};
test_label[279] = '{32'h4117e3b7};
test_output[279] = '{32'h429580dd};
/*############ DEBUG ############
test_input[2232:2239] = '{9.49309447474, -98.273201373, -81.446316435, 76.9828437765, -53.3666927817, -56.7037013664, -89.0805373018, 84.2440763371};
test_label[279] = '{9.49309447474};
test_output[279] = '{74.7516838579};
############ END DEBUG ############*/
test_input[2240:2247] = '{32'h421fb4ff, 32'h41af3754, 32'h3e34d87e, 32'hc1b6b5b9, 32'hbfa23247, 32'hc20a2f1d, 32'h428ae028, 32'h41a35bee};
test_label[280] = '{32'hc20a2f1d};
test_output[280] = '{32'h42cff7b6};
/*############ DEBUG ############
test_input[2240:2247] = '{39.9267541495, 21.9020155448, 0.176607105427, -22.8387314304, -1.26715932402, -34.5460080016, 69.4378039723, 20.4198870713};
test_label[280] = '{-34.5460080016};
test_output[280] = '{103.983811974};
############ END DEBUG ############*/
test_input[2248:2255] = '{32'h42886d4e, 32'hc1dee082, 32'h42b0d67b, 32'h4275ca29, 32'h424d687f, 32'h421258d1, 32'h42bf84fa, 32'hc15ffbba};
test_label[281] = '{32'h421258d1};
test_output[281] = '{32'h426cb1cd};
/*############ DEBUG ############
test_input[2248:2255] = '{68.2134864416, -27.8596238261, 88.4189077808, 61.447420233, 51.3520484134, 36.5867338725, 95.7597189417, -13.9989562628};
test_label[281] = '{36.5867338725};
test_output[281] = '{59.1736333832};
############ END DEBUG ############*/
test_input[2256:2263] = '{32'hc17e5ee8, 32'hc21ebe9f, 32'hc25891fd, 32'hc2c50b9a, 32'h422ea513, 32'h42bfce18, 32'hc24d60da, 32'hc2706199};
test_label[282] = '{32'hc21ebe9f};
test_output[282] = '{32'h430796b4};
/*############ DEBUG ############
test_input[2256:2263] = '{-15.8981701609, -39.6861528501, -54.142566601, -98.5226597131, 43.6612061936, 95.9025280171, -51.3445799779, -60.0953102042};
test_label[282] = '{-39.6861528501};
test_output[282] = '{135.588680867};
############ END DEBUG ############*/
test_input[2264:2271] = '{32'h4269048d, 32'h42109da2, 32'h42a50549, 32'h42ba7182, 32'h4217988a, 32'hc2b4cb60, 32'hc22603dd, 32'h4294eb38};
test_label[283] = '{32'h42a50549};
test_output[283] = '{32'h412b61da};
/*############ DEBUG ############
test_input[2264:2271] = '{58.2544460111, 36.1539372694, 82.5103245417, 93.2216920604, 37.898964638, -90.3972166249, -41.5037722427, 74.4594143117};
test_label[283] = '{82.5103245417};
test_output[283] = '{10.7113898157};
############ END DEBUG ############*/
test_input[2272:2279] = '{32'h42ba4da4, 32'hc28275dd, 32'h416af17e, 32'h4182a6a2, 32'h419e187d, 32'hc1ea0685, 32'h41ee3d8c, 32'hc25f6f8c};
test_label[284] = '{32'h419e187d};
test_output[284] = '{32'h4292c784};
/*############ DEBUG ############
test_input[2272:2279] = '{93.1516400451, -65.2302008303, 14.68395801, 16.3313642578, 19.7619577992, -29.2531840404, 29.7800516696, -55.8589343327};
test_label[284] = '{19.7619577992};
test_output[284] = '{73.3896822459};
############ END DEBUG ############*/
test_input[2280:2287] = '{32'h42b6029f, 32'hc28f8bad, 32'h42c78eae, 32'h419e9972, 32'hc2b8d047, 32'hc277c470, 32'hc203d277, 32'hc21053cb};
test_label[285] = '{32'hc277c470};
test_output[285] = '{32'h4321b87d};
/*############ DEBUG ############
test_input[2280:2287] = '{91.0051196817, -71.7728060551, 99.7786681096, 19.8249238936, -92.4067932229, -61.9418330454, -32.9555317766, -36.0818293983};
test_label[285] = '{-61.9418330454};
test_output[285] = '{161.720655916};
############ END DEBUG ############*/
test_input[2288:2295] = '{32'h42a5e378, 32'hc1f15118, 32'h423df6e1, 32'hc2a1b0fe, 32'h413d3c4a, 32'h4263ecd7, 32'h41b0fab6, 32'hc28046cb};
test_label[286] = '{32'h413d3c4a};
test_output[286] = '{32'h428e3bef};
/*############ DEBUG ############
test_input[2288:2295] = '{82.9442731934, -30.1645970167, 47.4910943846, -80.8456844702, 11.8272191209, 56.9812886174, 22.1224182123, -64.138266517};
test_label[286] = '{11.8272191209};
test_output[286] = '{71.1170540725};
############ END DEBUG ############*/
test_input[2296:2303] = '{32'h41ce2c87, 32'hc241a542, 32'h4289632e, 32'h3fa3e23d, 32'hc2030697, 32'hc2c1068e, 32'h42a26d3b, 32'h42bf42bd};
test_label[287] = '{32'hc241a542};
test_output[287] = '{32'h43100aaf};
/*############ DEBUG ############
test_input[2296:2303] = '{25.7717426488, -48.4113862083, 68.6937088544, 1.28034168544, -32.7564356028, -96.5128038021, 81.2133439151, 95.6303516143};
test_label[287] = '{-48.4113862083};
test_output[287] = '{144.041738371};
############ END DEBUG ############*/
test_input[2304:2311] = '{32'h3f356d43, 32'h41bf8bff, 32'h40153009, 32'hc1357da6, 32'hc259f6bf, 32'h42495b8b, 32'hc26bb79a, 32'hc0e6b097};
test_label[288] = '{32'hc0e6b097};
test_output[288] = '{32'h4266319d};
/*############ DEBUG ############
test_input[2304:2311] = '{0.708698456645, 23.9433570373, 2.33105677885, -11.3431762745, -54.4909635149, 50.3393957293, -58.9293000342, -7.20905623477};
test_label[288] = '{-7.20905623477};
test_output[288] = '{57.5484519641};
############ END DEBUG ############*/
test_input[2312:2319] = '{32'h4169d6c0, 32'h428ff2d8, 32'h425e9747, 32'hc1585171, 32'hc1afd2c5, 32'hc27e7ac0, 32'h40093b45, 32'hc28ef4df};
test_label[289] = '{32'hc28ef4df};
test_output[289] = '{32'h430f73dc};
/*############ DEBUG ############
test_input[2312:2319] = '{14.6149291281, 71.9743032727, 55.6477332825, -13.5198831438, -21.9779156776, -63.6198723814, 2.14424249065, -71.4782654936};
test_label[289] = '{-71.4782654936};
test_output[289] = '{143.452568848};
############ END DEBUG ############*/
test_input[2320:2327] = '{32'h42bbb6e6, 32'hc1826ecb, 32'h422b19af, 32'h42024c03, 32'h42827389, 32'hbfe94899, 32'h417fb90d, 32'hc1f59c32};
test_label[290] = '{32'h417fb90d};
test_output[290] = '{32'h429bbfc4};
/*############ DEBUG ############
test_input[2320:2327] = '{93.8572238041, -16.3040975364, 42.7750831423, 32.574231523, 65.2256526033, -1.82252796703, 15.982678723, -30.7012672643};
test_label[290] = '{15.982678723};
test_output[290] = '{77.8745450812};
############ END DEBUG ############*/
test_input[2328:2335] = '{32'h42ac96a1, 32'hc289567a, 32'h427920a6, 32'h4220aa6a, 32'h4252a3e5, 32'h429c6bfc, 32'h42b3d826, 32'hc22ad6b0};
test_label[291] = '{32'h42ac96a1};
test_output[291] = '{32'h4069de76};
/*############ DEBUG ############
test_input[2328:2335] = '{86.2941960851, -68.6689010981, 62.2818843363, 40.16642097, 52.6600540364, 78.2109051476, 89.9221679089, -42.7096546551};
test_label[291] = '{86.2941960851};
test_output[291] = '{3.65420297851};
############ END DEBUG ############*/
test_input[2336:2343] = '{32'hc29472bd, 32'h429f814d, 32'h4296aba9, 32'h42a71274, 32'hc1fba744, 32'h41777342, 32'h41ebddbf, 32'h41065ade};
test_label[292] = '{32'h42a71274};
test_output[292] = '{32'h3cba6be5};
/*############ DEBUG ############
test_input[2336:2343] = '{-74.2240973163, 79.7525416765, 75.3352770508, 83.5360401181, -31.4566725167, 15.4656387061, 29.4832750007, 8.39718400072};
test_label[292] = '{83.5360401181};
test_output[292] = '{0.0227565260659};
############ END DEBUG ############*/
test_input[2344:2351] = '{32'hc29ba60e, 32'hc24e98fb, 32'hc27f7c9b, 32'hc2915b1e, 32'hc23af587, 32'hc1095d11, 32'hc2ad498e, 32'hc20b8388};
test_label[293] = '{32'hc20b8388};
test_output[293] = '{32'h41d25887};
/*############ DEBUG ############
test_input[2344:2351] = '{-77.8243269495, -51.6493966788, -63.8716869028, -72.6779643124, -46.7397735938, -8.58522112387, -86.6436629255, -34.8784477613};
test_label[293] = '{-34.8784477613};
test_output[293] = '{26.2932266374};
############ END DEBUG ############*/
test_input[2352:2359] = '{32'h42c37f7e, 32'h4289050d, 32'hc2169069, 32'hc2066d34, 32'h42427ed7, 32'h4140a93f, 32'h42217f95, 32'h42281dba};
test_label[294] = '{32'h42c37f7e};
test_output[294] = '{32'h2a618000};
/*############ DEBUG ############
test_input[2352:2359] = '{97.7490073409, 68.5098647617, -37.6410253215, -33.6066443641, 48.6238664341, 12.041320079, 40.3745900879, 42.0290280691};
test_label[294] = '{97.7490073409};
test_output[294] = '{2.00284233642e-13};
############ END DEBUG ############*/
test_input[2360:2367] = '{32'h41d8d599, 32'h427ca96d, 32'h41a671a0, 32'h428b72d8, 32'h428222b6, 32'h4206ce64, 32'hc1dea523, 32'h42817ce9};
test_label[295] = '{32'hc1dea523};
test_output[295] = '{32'h42c32528};
/*############ DEBUG ############
test_input[2360:2367] = '{27.1042965465, 63.1654558951, 20.8054804904, 69.7243073783, 65.0677924954, 33.7015517506, -27.8306323449, 64.7439657346};
test_label[295] = '{-27.8306323449};
test_output[295] = '{97.5725720942};
############ END DEBUG ############*/
test_input[2368:2375] = '{32'hc206379f, 32'hc20070f1, 32'h426413db, 32'hc2b5074a, 32'hc2c1602a, 32'hc2b47219, 32'hc2a3428c, 32'h41e3c28c};
test_label[296] = '{32'h426413db};
test_output[296] = '{32'h2ae0b000};
/*############ DEBUG ############
test_input[2368:2375] = '{-33.5543164947, -32.1102932592, 57.0193882693, -90.5142374403, -96.6878211308, -90.2228464867, -81.6299778758, 28.4699931894};
test_label[296] = '{57.0193882693};
test_output[296] = '{3.99125177353e-13};
############ END DEBUG ############*/
test_input[2376:2383] = '{32'h42037e4b, 32'hc2488aee, 32'h41a003b4, 32'h4118f3bc, 32'hc1e32d54, 32'hc0946efd, 32'hc21f1f22, 32'hc2b66a4b};
test_label[297] = '{32'h4118f3bc};
test_output[297] = '{32'h41ba82b9};
/*############ DEBUG ############
test_input[2376:2383] = '{32.8733323975, -50.1356741224, 20.0018075976, 9.55950577489, -28.3971325723, -4.63854850929, -39.7804019757, -91.2076053258};
test_label[297] = '{9.55950577489};
test_output[297] = '{23.3138291929};
############ END DEBUG ############*/
test_input[2384:2391] = '{32'h4212009d, 32'h42b6c669, 32'hc1f60f85, 32'h420ee677, 32'hc277c82b, 32'hc2a009cd, 32'h42539e9b, 32'hc180726e};
test_label[298] = '{32'hc2a009cd};
test_output[298] = '{32'h432b681b};
/*############ DEBUG ############
test_input[2384:2391] = '{36.5005978358, 91.3875169323, -30.7575784664, 35.7250633294, -61.9454784165, -80.01914026, 52.9048864371, -16.0558731354};
test_label[298] = '{-80.01914026};
test_output[298] = '{171.406657192};
############ END DEBUG ############*/
test_input[2392:2399] = '{32'hc28b76bc, 32'hc2b8664d, 32'hc17cc02d, 32'hc2704c0c, 32'hc2446e8a, 32'h42bbb86e, 32'hc219018a, 32'hc258f4c4};
test_label[299] = '{32'hc17cc02d};
test_output[299] = '{32'h42db5073};
/*############ DEBUG ############
test_input[2392:2399] = '{-69.7319026163, -92.199807774, -15.796917699, -60.0742646798, -49.1079486567, 93.8602111846, -38.2515039215, -54.239029036};
test_label[299] = '{-15.796917699};
test_output[299] = '{109.657128884};
############ END DEBUG ############*/
test_input[2400:2407] = '{32'hc2086f67, 32'hc286fb3c, 32'h42003b15, 32'h41bf576c, 32'hc18ad48e, 32'hc2998116, 32'hc271b1f0, 32'h42800d6d};
test_label[300] = '{32'hc286fb3c};
test_output[300] = '{32'h43038455};
/*############ DEBUG ############
test_input[2400:2407] = '{-34.1087914466, -67.4906918429, 32.0576961619, 23.9176855521, -17.3537869364, -76.7521227384, -60.4237682139, 64.0262243024};
test_label[300] = '{-67.4906918429};
test_output[300] = '{131.516916145};
############ END DEBUG ############*/
test_input[2408:2415] = '{32'hc206f20a, 32'h42b2abf7, 32'h3fc8cab9, 32'hc1c19eea, 32'hc28ced0e, 32'hc07b3ef4, 32'hc184138d, 32'hc2c18a32};
test_label[301] = '{32'h3fc8cab9};
test_output[301] = '{32'h42af88cc};
/*############ DEBUG ############
test_input[2408:2415] = '{-33.7363669214, 89.3358714619, 1.56868662154, -24.2025953448, -70.4629961188, -3.92571725342, -16.5095471084, -96.7699119195};
test_label[301] = '{1.56868662154};
test_output[301] = '{87.7671848404};
############ END DEBUG ############*/
test_input[2416:2423] = '{32'h42156918, 32'h41b0db22, 32'h42469cde, 32'h40c64d1f, 32'hc26b72c8, 32'hc28b0d8d, 32'hc279c097, 32'hc204cec8};
test_label[302] = '{32'hc28b0d8d};
test_output[302] = '{32'h42ee5bfc};
/*############ DEBUG ############
test_input[2416:2423] = '{37.3526296915, 22.1069991272, 49.6531906404, 6.19691429539, -58.8620904051, -69.5264642083, -62.4380743172, -33.2019350672};
test_label[302] = '{-69.5264642083};
test_output[302] = '{119.179659398};
############ END DEBUG ############*/
test_input[2424:2431] = '{32'h418f6f37, 32'h4216e7d3, 32'hc2b50a3c, 32'hc2b64965, 32'hc2acf6ed, 32'h4288b080, 32'hc234555c, 32'hc0f3dafd};
test_label[303] = '{32'hc2acf6ed};
test_output[303] = '{32'h431ad3b7};
/*############ DEBUG ############
test_input[2424:2431] = '{17.9293046416, 37.7263926669, -90.519989588, -91.1433523639, -86.4822770796, 68.3447277775, -45.0833600819, -7.62048183025};
test_label[303] = '{-86.4822770796};
test_output[303] = '{154.827004857};
############ END DEBUG ############*/
test_input[2432:2439] = '{32'h3edbd253, 32'hc283800a, 32'hc1a99d99, 32'h425d0eeb, 32'hc1863792, 32'hc1c0a1f7, 32'h421905c0, 32'hc1442d0e};
test_label[304] = '{32'h421905c0};
test_output[304] = '{32'h41881255};
/*############ DEBUG ############
test_input[2432:2439] = '{0.429339030391, -65.7500737286, -21.2019516163, 55.2645681437, -16.7771341448, -24.0790837412, 38.2556163227, -12.2609993873};
test_label[304] = '{38.2556163227};
test_output[304] = '{17.0089518621};
############ END DEBUG ############*/
test_input[2440:2447] = '{32'h405e3ed3, 32'h4003b25f, 32'h41aef0d5, 32'hc2089014, 32'hc24694d2, 32'hc268973a, 32'h422c863c, 32'hc27a2fbf};
test_label[305] = '{32'h422c863c};
test_output[305] = '{32'h302025e2};
/*############ DEBUG ############
test_input[2440:2447] = '{3.47258440961, 2.05776179269, 21.8675947128, -34.1407014603, -49.6453320738, -58.1476828211, 43.1310894959, -62.5466275746};
test_label[305] = '{43.1310894959};
test_output[305] = '{5.82614956449e-10};
############ END DEBUG ############*/
test_input[2448:2455] = '{32'h429e9940, 32'h410b86c7, 32'h40bf5c2f, 32'hc28bd92e, 32'h4089cdd9, 32'hc119385d, 32'h3fc7a6e3, 32'h42c26c8f};
test_label[306] = '{32'h410b86c7};
test_output[306] = '{32'h42b0fbb6};
/*############ DEBUG ############
test_input[2448:2455] = '{79.2993131508, 8.72040472328, 5.9800027505, -69.9241778472, 4.30637809806, -9.57626039832, 1.55978045266, 97.2120285748};
test_label[306] = '{8.72040472328};
test_output[306] = '{88.4916238681};
############ END DEBUG ############*/
test_input[2456:2463] = '{32'hc2707d45, 32'h414c36d2, 32'h42bd5079, 32'hc164f699, 32'hc1210402, 32'hc1a623ba, 32'h42b36747, 32'h42303d1e};
test_label[307] = '{32'h42bd5079};
test_output[307] = '{32'h3be60927};
/*############ DEBUG ############
test_input[2456:2463] = '{-60.1223328289, 12.7633837165, 94.6571758002, -14.3102049523, -10.0634786683, -20.7674439052, 89.7017149392, 44.0596838334};
test_label[307] = '{94.6571758002};
test_output[307] = '{0.00702013393999};
############ END DEBUG ############*/
test_input[2464:2471] = '{32'h42252dfc, 32'h42b45850, 32'h42169551, 32'hc2811d35, 32'h429e6817, 32'hc2b51720, 32'hc29d3241, 32'hc190c966};
test_label[308] = '{32'hc2b51720};
test_output[308] = '{32'h4334b7b9};
/*############ DEBUG ############
test_input[2464:2471] = '{41.2949054106, 90.172485827, 37.6458184079, -64.5570432875, 79.2033031957, -90.5451684466, -78.5981502801, -18.0983395941};
test_label[308] = '{-90.5451684466};
test_output[308] = '{180.717671498};
############ END DEBUG ############*/
test_input[2472:2479] = '{32'hc22ebc26, 32'hc283f701, 32'hc2345c45, 32'hc2192e7b, 32'hc25f2e10, 32'h42c27b45, 32'h423a164f, 32'hc2b5939e};
test_label[309] = '{32'h423a164f};
test_output[309] = '{32'h424ae03b};
/*############ DEBUG ############
test_input[2472:2479] = '{-43.6837387242, -65.9824281018, -45.0901071961, -38.2953903721, -55.7949816575, 97.2407577916, 46.5217840434, -90.7883155374};
test_label[309] = '{46.5217840434};
test_output[309] = '{50.7189737482};
############ END DEBUG ############*/
test_input[2480:2487] = '{32'h424ca0d0, 32'hc20d4d2c, 32'hc18e84e5, 32'h41d2a363, 32'hc1bd132e, 32'hc25bb8d9, 32'h429de756, 32'h42011959};
test_label[310] = '{32'h41d2a363};
test_output[310] = '{32'h42527cfb};
/*############ DEBUG ############
test_input[2480:2487] = '{51.157045302, -35.325361753, -17.8148890751, 26.3297795474, -23.6343646902, -54.9305151446, 78.95182978, 32.2747530923};
test_label[310] = '{26.3297795474};
test_output[310] = '{52.6220502326};
############ END DEBUG ############*/
test_input[2488:2495] = '{32'h42aa08a0, 32'h4174ba5b, 32'h41d9f9a0, 32'h4297dc58, 32'h429edbd8, 32'hc2486433, 32'hc230f7f7, 32'h412ebb4c};
test_label[311] = '{32'h4297dc58};
test_output[311] = '{32'h41117203};
/*############ DEBUG ############
test_input[2488:2495] = '{85.016844797, 15.2954970616, 27.2468870042, 75.9303604443, 79.4293834962, -50.0978525445, -44.2421541189, 10.9207267158};
test_label[311] = '{75.9303604443};
test_output[311] = '{9.09033463821};
############ END DEBUG ############*/
test_input[2496:2503] = '{32'h420fefec, 32'h4246e200, 32'hc2c25e4f, 32'h4281e9bb, 32'hc2ac81d4, 32'h42068226, 32'hc29ae069, 32'h4266b9b5};
test_label[312] = '{32'h4246e200};
test_output[312] = '{32'h4173c8b1};
/*############ DEBUG ############
test_input[2496:2503] = '{35.9842992574, 49.720701478, -97.1841979368, 64.9565056256, -86.2535672564, 33.6270971288, -77.4383026309, 57.6813557206};
test_label[312] = '{49.720701478};
test_output[312] = '{15.2364966857};
############ END DEBUG ############*/
test_input[2504:2511] = '{32'hc20981b8, 32'h42111a7e, 32'hc2abdce7, 32'h428b62c7, 32'h40a561bf, 32'hc0d09ec8, 32'h42a3b658, 32'h415fd2bb};
test_label[313] = '{32'h40a561bf};
test_output[313] = '{32'h4299603d};
/*############ DEBUG ############
test_input[2504:2511] = '{-34.376677908, 36.275870566, -85.9314469913, 69.6929265249, 5.16818175551, -6.51938247307, 81.8561404507, 13.9889474461};
test_label[313] = '{5.16818175551};
test_output[313] = '{76.6879639141};
############ END DEBUG ############*/
test_input[2512:2519] = '{32'h42bc5f90, 32'h411d8241, 32'h416e5596, 32'hc29074ae, 32'h422b3cc9, 32'hc1260ebc, 32'h4293988e, 32'h41e0e446};
test_label[314] = '{32'h422b3cc9};
test_output[314] = '{32'h424d8258};
/*############ DEBUG ############
test_input[2512:2519] = '{94.1866479145, 9.84430064937, 14.8958948003, -72.2278866905, 42.8093599077, -10.3785970153, 73.7979595699, 28.1114617681};
test_label[314] = '{42.8093599077};
test_output[314] = '{51.3772880082};
############ END DEBUG ############*/
test_input[2520:2527] = '{32'hc2aa19ff, 32'hc1ec8085, 32'hc0c8a530, 32'hc287cff5, 32'hc1413d43, 32'h4292e3ec, 32'h425d6d83, 32'h429249a6};
test_label[315] = '{32'hc1413d43};
test_output[315] = '{32'h42ac2720};
/*############ DEBUG ############
test_input[2520:2527] = '{-85.0507767462, -29.5627543286, -6.27016460495, -67.9061634297, -12.0774568474, 73.4451633066, 55.3569432661, 73.1438427497};
test_label[315] = '{-12.0774568474};
test_output[315] = '{86.0764136467};
############ END DEBUG ############*/
test_input[2528:2535] = '{32'hc2b70986, 32'hc1be52dc, 32'hc22ee83a, 32'h42b6c0f9, 32'hc20601ea, 32'hbf2fc8fe, 32'hc2305d87, 32'hc25d160e};
test_label[316] = '{32'hbf2fc8fe};
test_output[316] = '{32'h42b8208b};
/*############ DEBUG ############
test_input[2528:2535] = '{-91.5186011808, -23.790459454, -43.7267835987, 91.3768985676, -33.5018679091, -0.686660650877, -44.0913357898, -55.2715375135};
test_label[316] = '{-0.686660650877};
test_output[316] = '{92.0635592185};
############ END DEBUG ############*/
test_input[2536:2543] = '{32'h428d2324, 32'h429e70c3, 32'hc2856ebc, 32'hc2b095d0, 32'h408dd2aa, 32'hc24a8d97, 32'h410077bc, 32'h42bdc9a8};
test_label[317] = '{32'hc24a8d97};
test_output[317] = '{32'h4311883a};
/*############ DEBUG ############
test_input[2536:2543] = '{70.568632981, 79.2202400053, -66.7162750594, -88.2926016905, 4.4319657023, -50.6382698605, 8.02923209384, 94.8938635506};
test_label[317] = '{-50.6382698605};
test_output[317] = '{145.532133567};
############ END DEBUG ############*/
test_input[2544:2551] = '{32'h42b00eb5, 32'hc1f9c61d, 32'h41c504a7, 32'hc2ba6586, 32'h429c8772, 32'hc1281672, 32'hc0ade969, 32'hc155e516};
test_label[318] = '{32'h41c504a7};
test_output[318] = '{32'h427d9b25};
/*############ DEBUG ############
test_input[2544:2551] = '{88.0287235298, -31.2217357767, 24.6272714743, -93.1982875338, 78.2645448688, -10.5054802313, -5.43474246578, -13.3684294267};
test_label[318] = '{24.6272714743};
test_output[318] = '{63.4015095278};
############ END DEBUG ############*/
test_input[2552:2559] = '{32'h42b9858e, 32'hc2bba61d, 32'h424020cc, 32'hc2b986f1, 32'h420965b8, 32'hc245d3ef, 32'hc219cfb1, 32'h4288a020};
test_label[319] = '{32'h4288a020};
test_output[319] = '{32'h41c395b7};
/*############ DEBUG ############
test_input[2552:2559] = '{92.7608470973, -93.8244384606, 48.0320266245, -92.763557152, 34.3493343232, -49.4569676396, -38.4528224328, 68.3127437299};
test_label[319] = '{68.3127437299};
test_output[319] = '{24.4481033675};
############ END DEBUG ############*/
test_input[2560:2567] = '{32'hc29d9bd1, 32'hc1b33234, 32'hc26bf204, 32'h42291c0c, 32'h425e4ea2, 32'hc20bac7e, 32'h40587f6c, 32'h42be7834};
test_label[320] = '{32'h40587f6c};
test_output[320] = '{32'h42b7b439};
/*############ DEBUG ############
test_input[2560:2567] = '{-78.8043321126, -22.3995136648, -58.9863449659, 42.277388842, 55.5767882448, -34.9184486181, 3.38277722426, 95.2347741316};
test_label[320] = '{3.38277722426};
test_output[320] = '{91.8519969073};
############ END DEBUG ############*/
test_input[2568:2575] = '{32'hc081f69e, 32'h428e4925, 32'h3f9a8ceb, 32'hc26a0989, 32'hc245626a, 32'hc2378c1f, 32'hc187dd2b, 32'hbf84c8d3};
test_label[321] = '{32'h428e4925};
test_output[321] = '{32'h80000000};
/*############ DEBUG ############
test_input[2568:2575] = '{-4.06135460591, 71.1428632319, 1.20742546685, -58.5093120923, -49.3461093052, -45.8868379845, -16.982991459, -1.03737863792};
test_label[321] = '{71.1428632319};
test_output[321] = '{-0.0};
############ END DEBUG ############*/
test_input[2576:2583] = '{32'hc25513b1, 32'hc26646c3, 32'hc28343db, 32'hc2920528, 32'h4261a15a, 32'hc273e30d, 32'hc2c73a86, 32'h42564587};
test_label[322] = '{32'h4261a15a};
test_output[322] = '{32'h3d68a7e7};
/*############ DEBUG ############
test_input[2576:2583] = '{-53.2692292429, -57.5691047873, -65.6325273241, -73.0100726668, 56.407570479, -60.971729937, -99.6143038731, 53.5678995232};
test_label[322] = '{56.407570479};
test_output[322] = '{0.0568007495389};
############ END DEBUG ############*/
test_input[2584:2591] = '{32'h424d1ca4, 32'h41c01716, 32'h41e599b5, 32'h4286410d, 32'h42b7cdb4, 32'h423a0542, 32'hc1bb9625, 32'h42c7015c};
test_label[323] = '{32'h41c01716};
test_output[323] = '{32'h4296fbd9};
/*############ DEBUG ############
test_input[2584:2591] = '{51.2779705806, 24.0112716311, 28.7000530317, 67.1270518154, 91.9017650181, 46.505136359, -23.4483118075, 99.502658699};
test_label[323] = '{24.0112716311};
test_output[323] = '{75.4918869474};
############ END DEBUG ############*/
test_input[2592:2599] = '{32'hc2aa46ca, 32'h423f385f, 32'h426d2862, 32'h4232855e, 32'hc236bbf3, 32'h40c2e46a, 32'h42c7ef90, 32'hc201b0b7};
test_label[324] = '{32'hc236bbf3};
test_output[324] = '{32'h4311a6c5};
/*############ DEBUG ############
test_input[2592:2599] = '{-85.1382580639, 47.8050511508, 59.2894358406, 44.6302396953, -45.6835452847, 6.09038243049, 99.9678958354, -32.422573028};
test_label[324] = '{-45.6835452847};
test_output[324] = '{145.65144112};
############ END DEBUG ############*/
test_input[2600:2607] = '{32'hc223ab08, 32'hc1f6ad44, 32'hc0b5d4f6, 32'h42873f75, 32'hc2586b79, 32'h419405ba, 32'h4299f72b, 32'h3f328ea5};
test_label[325] = '{32'hc223ab08};
test_output[325] = '{32'h42ebccba};
/*############ DEBUG ############
test_input[2600:2607] = '{-40.917021953, -30.8346025307, -5.68224614726, 67.6239360071, -54.1049522898, 18.5027963746, 76.9827518281, 0.697489104821};
test_label[325] = '{-40.917021953};
test_output[325] = '{117.89985998};
############ END DEBUG ############*/
test_input[2608:2615] = '{32'hc2af4a76, 32'hc244de5e, 32'hbffc91c1, 32'h42c77c90, 32'h426f43c8, 32'h41fe8fc8, 32'hc1f34ed0, 32'h423d8287};
test_label[326] = '{32'hbffc91c1};
test_output[326] = '{32'h42cb6ed7};
/*############ DEBUG ############
test_input[2608:2615] = '{-87.6454308543, -49.2171568363, -1.97319810385, 99.7432851147, 59.8161930413, 31.8202056898, -30.4134832035, 47.3774665923};
test_label[326] = '{-1.97319810385};
test_output[326] = '{101.716483219};
############ END DEBUG ############*/
test_input[2616:2623] = '{32'h41d648f3, 32'h4284db21, 32'hc1e085f2, 32'h4222fa10, 32'h41924556, 32'h41f10708, 32'h42171515, 32'hc2158ae9};
test_label[327] = '{32'h41d648f3};
test_output[327] = '{32'h421e91c9};
/*############ DEBUG ############
test_input[2616:2623] = '{26.7856206798, 66.4279886449, -28.0654027797, 40.7442022581, 18.2838551451, 30.128433251, 37.7705882465, -37.385654684};
test_label[327] = '{26.7856206798};
test_output[327] = '{39.6423679651};
############ END DEBUG ############*/
test_input[2624:2631] = '{32'h42aece14, 32'h42290650, 32'hc2af9478, 32'hc2b4f113, 32'hc2bae1ae, 32'h42c4b4c1, 32'hc28e1307, 32'hc2afa4cb};
test_label[328] = '{32'hc2afa4cb};
test_output[328] = '{32'h433a2cc7};
/*############ DEBUG ############
test_input[2624:2631] = '{87.4024948862, 42.2561634871, -87.7899805534, -90.4708489925, -93.4407804074, 98.3530332805, -71.0371662016, -87.8218606827};
test_label[328] = '{-87.8218606827};
test_output[328] = '{186.174911512};
############ END DEBUG ############*/
test_input[2632:2639] = '{32'hc2979a21, 32'h41d7da90, 32'h427eb09a, 32'h40d6f248, 32'h42959185, 32'h3fdfd0c8, 32'h419b67a2, 32'hc23bd97d};
test_label[329] = '{32'h41d7da90};
test_output[329] = '{32'h423f35c5};
/*############ DEBUG ############
test_input[2632:2639] = '{-75.8010332183, 26.9817201604, 63.6724621236, 6.71707511754, 74.7842162792, 1.7485589551, 19.4256024022, -46.9623918986};
test_label[329] = '{26.9817201604};
test_output[329] = '{47.8025110545};
############ END DEBUG ############*/
test_input[2640:2647] = '{32'h42880e99, 32'h421990ca, 32'hc1d7901c, 32'hc24269eb, 32'h421a48eb, 32'hc2674984, 32'h42bc174c, 32'h42a49916};
test_label[330] = '{32'hc24269eb};
test_output[330] = '{32'h430ea621};
/*############ DEBUG ############
test_input[2640:2647] = '{68.0285104542, 38.3913946181, -26.9453663546, -48.6034355031, 38.5712097275, -57.8217928713, 94.0455035204, 82.2989941167};
test_label[330] = '{-48.6034355031};
test_output[330] = '{142.64894694};
############ END DEBUG ############*/
test_input[2648:2655] = '{32'h4294c23b, 32'hc293a974, 32'h428b8aad, 32'hc1ef1abd, 32'hc2c7bcd2, 32'h4162ae5b, 32'h41e30e48, 32'h415d888a};
test_label[331] = '{32'hc2c7bcd2};
test_output[331] = '{32'h432e4210};
/*############ DEBUG ############
test_input[2648:2655] = '{74.3793565059, -73.8309595512, 69.770849829, -29.8880549457, -99.8687873419, 14.1675672582, 28.3819742012, 13.8458347698};
test_label[331] = '{-99.8687873419};
test_output[331] = '{174.258061199};
############ END DEBUG ############*/
test_input[2656:2663] = '{32'hc15b68d3, 32'hc29c4610, 32'hc2074b4a, 32'hc1a0d6a2, 32'hc299f6e9, 32'hc29d88d7, 32'hc120ad44, 32'hc2546baf};
test_label[332] = '{32'hc2074b4a};
test_output[332] = '{32'h41be7383};
/*############ DEBUG ############
test_input[2656:2663] = '{-13.7130919142, -78.1368405383, -33.8235246316, -20.1048013559, -76.9822461263, -78.7672679056, -10.042300877, -53.1051614708};
test_label[332] = '{-33.8235246316};
test_output[332] = '{23.806403053};
############ END DEBUG ############*/
test_input[2664:2671] = '{32'hc2c29670, 32'h421d5468, 32'hc1d1b7cc, 32'hc192c6f7, 32'hc26a6ee9, 32'h42519f84, 32'hc13ae9dc, 32'hc1ac77fd};
test_label[333] = '{32'h42519f84};
test_output[333] = '{32'h360cf5b7};
/*############ DEBUG ############
test_input[2664:2671] = '{-97.2938246665, 39.3324276996, -26.2147438262, -18.3471513215, -58.6083088212, 52.4057784005, -11.6820949412, -21.5585874719};
test_label[333] = '{52.4057784005};
test_output[333] = '{2.10046512202e-06};
############ END DEBUG ############*/
test_input[2672:2679] = '{32'h41ff5da3, 32'h42570668, 32'h4168ca4e, 32'h41d7945d, 32'h41e67deb, 32'h4297938c, 32'hc2005214, 32'hc0f4bb70};
test_label[334] = '{32'h41d7945d};
test_output[334] = '{32'h42435ce9};
/*############ DEBUG ############
test_input[2672:2679] = '{31.9207201272, 53.7562578668, 14.5493908119, 26.9474439493, 28.8114836204, 75.7881781708, -32.0801543573, -7.64788062559};
test_label[334] = '{26.9474439493};
test_output[334] = '{48.8407342218};
############ END DEBUG ############*/
test_input[2680:2687] = '{32'h4207a87a, 32'hc290eb3a, 32'h41578896, 32'h415640d9, 32'hc210521a, 32'hc10a6d28, 32'hc2bcacea, 32'h418e9598};
test_label[335] = '{32'h418e9598};
test_output[335] = '{32'h4180bb5b};
/*############ DEBUG ############
test_input[2680:2687] = '{33.9145263483, -72.4594295089, 13.4708458627, 13.3908320101, -36.0801765426, -8.65164963802, -94.3377227985, 17.8230445372};
test_label[335] = '{17.8230445372};
test_output[335] = '{16.0914819164};
############ END DEBUG ############*/
test_input[2688:2695] = '{32'hc2896f00, 32'h429d69e1, 32'hc2bec3a0, 32'hc03c1090, 32'hbf7fd92d, 32'h42bbaf7e, 32'hc2890953, 32'hc2bfa66a};
test_label[336] = '{32'hc2896f00};
test_output[336] = '{32'h43228f3f};
/*############ DEBUG ############
test_input[2688:2695] = '{-68.7167978988, 78.7067942592, -95.3820799228, -2.93851083479, -0.999407594039, 93.8427556159, -68.5182145868, -95.8250274167};
test_label[336] = '{-68.7167978988};
test_output[336] = '{162.559553782};
############ END DEBUG ############*/
test_input[2696:2703] = '{32'h422457f6, 32'h42914b0e, 32'h417d25e8, 32'hc1923088, 32'hc2a17662, 32'hc2687493, 32'hc10e231e, 32'hc1bac932};
test_label[337] = '{32'hc1bac932};
test_output[337] = '{32'h42bffd5a};
/*############ DEBUG ############
test_input[2696:2703] = '{41.0859002091, 72.6465883869, 15.8217543788, -18.2736963, -80.7312175459, -58.1138404308, -8.88357399931, -23.3482402125};
test_label[337] = '{-23.3482402125};
test_output[337] = '{95.9948285994};
############ END DEBUG ############*/
test_input[2704:2711] = '{32'h424b25a7, 32'hc12de30e, 32'hc1553ab8, 32'h427c88d3, 32'hc13dbffb, 32'hc2374a89, 32'h4060e870, 32'h42bac6a3};
test_label[338] = '{32'h42bac6a3};
test_output[338] = '{32'h29a34000};
/*############ DEBUG ############
test_input[2704:2711] = '{50.786771323, -10.8679331783, -13.3268359825, 63.1336165501, -11.8593706741, -45.822787477, 3.51418682188, 93.3879637574};
test_label[338] = '{93.3879637574};
test_output[338] = '{7.2497563508e-14};
############ END DEBUG ############*/
test_input[2712:2719] = '{32'h42703afe, 32'h40ad73f8, 32'hc25e6047, 32'hc1939df3, 32'h429d66b3, 32'h40d20a02, 32'hc2c14300, 32'h4098479e};
test_label[339] = '{32'h4098479e};
test_output[339] = '{32'h4293e239};
/*############ DEBUG ############
test_input[2712:2719] = '{60.0576076705, 5.42040646929, -55.594020524, -18.4521245836, 78.7005821203, 6.56372169192, -96.630859231, 4.75874244807};
test_label[339] = '{4.75874244807};
test_output[339] = '{73.9418396802};
############ END DEBUG ############*/
test_input[2720:2727] = '{32'hc1a3de7b, 32'hc248be96, 32'hc21f6928, 32'hc18e39a7, 32'hc2613d84, 32'h42c51399, 32'hc18f2e62, 32'h41574e2b};
test_label[340] = '{32'hc18e39a7};
test_output[340] = '{32'h42e8a203};
/*############ DEBUG ############
test_input[2720:2727] = '{-20.4836338256, -50.1861194998, -39.8526933797, -17.7781499831, -56.3100729608, 98.5382773734, -17.8976473775, 13.4565836424};
test_label[340] = '{-17.7781499831};
test_output[340] = '{116.316427357};
############ END DEBUG ############*/
test_input[2728:2735] = '{32'hc2822f45, 32'h42b28db8, 32'hc2c6c7c0, 32'h419e18ef, 32'hc28658cd, 32'h424ae070, 32'h4226870a, 32'h422327f5};
test_label[341] = '{32'h419e18ef};
test_output[341] = '{32'h428b077c};
/*############ DEBUG ############
test_input[2728:2735] = '{-65.0923217129, 89.2767913335, -99.3901350847, 19.7621746973, -67.1734354084, 50.7191770963, 41.6318759233, 40.7890190737};
test_label[341] = '{19.7621746973};
test_output[341] = '{69.5146166362};
############ END DEBUG ############*/
test_input[2736:2743] = '{32'hc291f3f5, 32'h413c3e84, 32'hc2ad8a69, 32'hc23c0ab6, 32'hc05f7cfa, 32'hc288d4cf, 32'h4164811e, 32'h42b29162};
test_label[342] = '{32'hc288d4cf};
test_output[342] = '{32'h431db318};
/*############ DEBUG ############
test_input[2736:2743] = '{-72.9764775307, 11.765262487, -86.7703359927, -47.0104601022, -3.49200303004, -68.4156393106, 14.2815225633, 89.2839494087};
test_label[342] = '{-68.4156393106};
test_output[342] = '{157.699588719};
############ END DEBUG ############*/
test_input[2744:2751] = '{32'hc286c793, 32'h4296b73f, 32'h42b816f8, 32'h40a2a8c2, 32'hc20249f4, 32'h42c37831, 32'h42a63bd2, 32'hc28062c6};
test_label[343] = '{32'h42b816f8};
test_output[343] = '{32'h40b62f2f};
/*############ DEBUG ############
test_input[2744:2751] = '{-67.3897939719, 75.3578999463, 92.0448608801, 5.08310052277, -32.5722182743, 97.7347458234, 83.1168386029, -64.1929199324};
test_label[343] = '{92.0448608801};
test_output[343] = '{5.69325967275};
############ END DEBUG ############*/
test_input[2752:2759] = '{32'h424aed28, 32'hc2172d2d, 32'hc21da321, 32'hc16f0857, 32'hc0471db2, 32'hc2430c6d, 32'h421ada3b, 32'hc281a8b8};
test_label[344] = '{32'hc21da321};
test_output[344] = '{32'h42b44825};
/*############ DEBUG ############
test_input[2752:2759] = '{50.7315986561, -37.7941164829, -39.4093061538, -14.9395363201, -3.11118747495, -48.7621327113, 38.7131156607, -64.8295292038};
test_label[344] = '{-39.4093061538};
test_output[344] = '{90.1409108416};
############ END DEBUG ############*/
test_input[2760:2767] = '{32'h41fe992a, 32'hc21d8a40, 32'hc1d3e8da, 32'h41c04b55, 32'h41c74e5c, 32'h42a88f2e, 32'hc13f0f82, 32'h409661c7};
test_label[345] = '{32'h409661c7};
test_output[345] = '{32'h429f2912};
/*############ DEBUG ############
test_input[2760:2767] = '{31.8247880556, -39.385009871, -26.4886967165, 24.0367832072, 24.9132621446, 84.2796474684, -11.9412862028, 4.6994357969};
test_label[345] = '{4.6994357969};
test_output[345] = '{79.5802116715};
############ END DEBUG ############*/
test_input[2768:2775] = '{32'hc29d8c86, 32'hc29eb4a0, 32'h424ad84b, 32'h41c0ac7c, 32'h41bea428, 32'hc1859a59, 32'hc284db77, 32'hc2a95225};
test_label[346] = '{32'hc1859a59};
test_output[346] = '{32'h4286d2bc};
/*############ DEBUG ############
test_input[2768:2775] = '{-78.7744595037, -79.3527857814, 50.7112238099, 24.0842210587, 23.8301535812, -16.7003649681, -66.4286385906, -84.6604373471};
test_label[346] = '{-16.7003649681};
test_output[346] = '{67.411588778};
############ END DEBUG ############*/
test_input[2776:2783] = '{32'h4182648c, 32'hc212b3ac, 32'hc1faa31a, 32'h42a79de3, 32'h4239ae45, 32'h423168fc, 32'hc28e5e74, 32'hc1fc09e6};
test_label[347] = '{32'h4182648c};
test_output[347] = '{32'h428704c0};
/*############ DEBUG ############
test_input[2776:2783] = '{16.299094644, -36.6754625207, -31.3296399286, 83.8083716944, 46.4201833392, 44.3525228335, -71.1844756341, -31.5048333208};
test_label[347] = '{16.299094644};
test_output[347] = '{67.5092770504};
############ END DEBUG ############*/
test_input[2784:2791] = '{32'hc24952be, 32'h418e4b4d, 32'h42134aac, 32'hc267e3ed, 32'hc217e676, 32'h4240f02f, 32'hc1a2f808, 32'h401fc5b8};
test_label[348] = '{32'h401fc5b8};
test_output[348] = '{32'h4236f3d7};
/*############ DEBUG ############
test_input[2784:2791] = '{-50.3308010999, 17.7867678645, 36.8229206634, -57.9725834719, -37.9750581559, 48.2345560851, -20.3711098208, 2.49644274252};
test_label[348] = '{2.49644274252};
test_output[348] = '{45.7381244085};
############ END DEBUG ############*/
test_input[2792:2799] = '{32'hc23db206, 32'hc2379088, 32'h427706fa, 32'h429bb32e, 32'h411b5323, 32'h423397b6, 32'hc1ca6d8a, 32'hc26c743e};
test_label[349] = '{32'h427706fa};
test_output[349] = '{32'h4180bec2};
/*############ DEBUG ############
test_input[2792:2799] = '{-47.4238521415, -45.8911454477, 61.7568137414, 77.8499566559, 9.70779731218, 44.8981537094, -25.3034864312, -59.1135172764};
test_label[349] = '{61.7568137414};
test_output[349] = '{16.0931430169};
############ END DEBUG ############*/
test_input[2800:2807] = '{32'hc0ae5577, 32'h41a350de, 32'h4216c0f3, 32'hc22e7273, 32'hc2a26ac8, 32'h42ae2869, 32'hc212ffbf, 32'h41e07ee3};
test_label[350] = '{32'h4216c0f3};
test_output[350] = '{32'h42458fdf};
/*############ DEBUG ############
test_input[2800:2807] = '{-5.44793251112, 20.4144855888, 37.6884287445, -43.611765161, -81.2085575448, 87.0789267552, -36.7497518439, 28.0619570654};
test_label[350] = '{37.6884287445};
test_output[350] = '{49.3904980107};
############ END DEBUG ############*/
test_input[2808:2815] = '{32'hc0caebd2, 32'hc28ca948, 32'h4293055b, 32'hc2250082, 32'h41876bc5, 32'h42318032, 32'hc1fc88b5, 32'h420e5202};
test_label[351] = '{32'hc2250082};
test_output[351] = '{32'h42e5859c};
/*############ DEBUG ############
test_input[2808:2815] = '{-6.34128653713, -70.3306260558, 73.510462334, -41.2504948199, 16.9276220978, 44.3751891737, -31.5667520584, 35.5800873144};
test_label[351] = '{-41.2504948199};
test_output[351] = '{114.760957154};
############ END DEBUG ############*/
test_input[2816:2823] = '{32'h4055eb4d, 32'hc17b85e1, 32'h41b521f6, 32'hc13c8bc1, 32'hc29651d2, 32'hc29892d2, 32'h42a27f9f, 32'h411632e6};
test_label[352] = '{32'hc29651d2};
test_output[352] = '{32'h431c68b8};
/*############ DEBUG ############
test_input[2816:2823] = '{3.3424865842, -15.7201850101, 22.641581753, -11.7841193238, -75.1598019614, -76.2867566105, 81.249258945, 9.38742677164};
test_label[352] = '{-75.1598019614};
test_output[352] = '{156.409060906};
############ END DEBUG ############*/
test_input[2824:2831] = '{32'h426767da, 32'h4170c08f, 32'hc21cacd0, 32'hc1f6be96, 32'hc190c802, 32'hc287d076, 32'hc2a6fab3, 32'h4240d234};
test_label[353] = '{32'hc1f6be96};
test_output[353] = '{32'h42b1639b};
/*############ DEBUG ############
test_input[2824:2831] = '{57.8514183603, 15.0470118294, -39.1687619989, -30.8430596944, -18.0976599846, -67.9071531173, -83.4896479509, 48.2052781218};
test_label[353] = '{-30.8430596944};
test_output[353] = '{88.6945427273};
############ END DEBUG ############*/
test_input[2832:2839] = '{32'hc238f48c, 32'hc29bdbf1, 32'hc1f90434, 32'h423efac3, 32'h4270cff7, 32'h4200a4c9, 32'h41868d76, 32'hc253b1f1};
test_label[354] = '{32'h423efac3};
test_output[354] = '{32'h414754d4};
/*############ DEBUG ############
test_input[2832:2839] = '{-46.2388153101, -77.9295763637, -31.1270529583, 47.7448856674, 60.2030920514, 32.1609234429, 16.8190735062, -52.9237705055};
test_label[354] = '{47.7448856674};
test_output[354] = '{12.4582102696};
############ END DEBUG ############*/
test_input[2840:2847] = '{32'h41de30b5, 32'h419089bf, 32'hc0f706f1, 32'h425feed3, 32'h41bb4dde, 32'hc299218c, 32'h42a1989a, 32'h418c8bc2};
test_label[355] = '{32'h419089bf};
test_output[355] = '{32'h427aec56};
/*############ DEBUG ############
test_input[2840:2847] = '{27.7737836648, 18.0672585128, -7.71959727118, 55.9832249803, 23.413020623, -76.5655229491, 80.7980535199, 17.5682418222};
test_label[355] = '{18.0672585128};
test_output[355] = '{62.7307950072};
############ END DEBUG ############*/
test_input[2848:2855] = '{32'hc28c3b62, 32'h425f1b9b, 32'h413b0155, 32'h42881928, 32'hc28843a5, 32'h4252bb3b, 32'hc2513a93, 32'h428ff571};
test_label[356] = '{32'h4252bb3b};
test_output[356] = '{32'h419a8722};
/*############ DEBUG ############
test_input[2848:2855] = '{-70.1159852363, 55.7769568712, 11.6878251624, 68.0491342, -68.1321210745, 52.6828413461, -52.307200278, 71.9793763039};
test_label[356] = '{52.6828413461};
test_output[356] = '{19.315983614};
############ END DEBUG ############*/
test_input[2856:2863] = '{32'h42a5d62c, 32'hc252bc98, 32'hc1fcc080, 32'hc1c8a547, 32'hc29683eb, 32'h40aef63c, 32'h421eb4e1, 32'hc1ebf8b7};
test_label[357] = '{32'hc1ebf8b7};
test_output[357] = '{32'h42e0d45a};
/*############ DEBUG ############
test_input[2856:2863] = '{82.9183019665, -52.6841737357, -31.5939938957, -25.0807010122, -75.2576512021, 5.46755792758, 39.6766406981, -29.496443437};
test_label[357] = '{-29.496443437};
test_output[357] = '{112.414745403};
############ END DEBUG ############*/
test_input[2864:2871] = '{32'h42b4d410, 32'h42bb65cd, 32'hc24688c0, 32'hc229aca7, 32'h412e90c6, 32'h42c21600, 32'hc12f497d, 32'h41fe6bf4};
test_label[358] = '{32'h42bb65cd};
test_output[358] = '{32'h40585375};
/*############ DEBUG ############
test_input[2864:2871] = '{90.4141816459, 93.6988331183, -49.6335457223, -42.4186066783, 10.910344966, 97.0429688181, -10.9554418846, 31.8027116149};
test_label[358] = '{93.6988331183};
test_output[358] = '{3.38009385522};
############ END DEBUG ############*/
test_input[2872:2879] = '{32'hc1d50a7b, 32'h41c46681, 32'hc096a892, 32'h42c0e39b, 32'hc23ef818, 32'h40bdb905, 32'h428913e4, 32'h42478479};
test_label[359] = '{32'h428913e4};
test_output[359] = '{32'h41df3edb};
/*############ DEBUG ############
test_input[2872:2879] = '{-26.6301175861, 24.5500507858, -4.70807748589, 96.4445434972, -47.7422775178, 5.92883559375, 68.5388523946, 49.8793693213};
test_label[359] = '{68.5388523946};
test_output[359] = '{27.9056911026};
############ END DEBUG ############*/
test_input[2880:2887] = '{32'hc2310703, 32'hc2826e5d, 32'h41625a0b, 32'h42441644, 32'hc0fcc375, 32'h41b9dd73, 32'h42266e36, 32'h423c13f1};
test_label[360] = '{32'h42266e36};
test_output[360] = '{32'h40f15262};
/*############ DEBUG ############
test_input[2880:2887] = '{-44.2568467707, -65.2155555213, 14.1469830722, 49.0217451871, -7.89885970169, 23.2331293264, 41.6076271994, 47.0194752974};
test_label[360] = '{41.6076271994};
test_output[360] = '{7.54130653623};
############ END DEBUG ############*/
test_input[2888:2895] = '{32'h425928cd, 32'h42a48bee, 32'hc29b9d55, 32'h41a037a4, 32'h42997d17, 32'hc204909e, 32'hc29d9a80, 32'hc20be98a};
test_label[361] = '{32'h41a037a4};
test_output[361] = '{32'h42790019};
/*############ DEBUG ############
test_input[2888:2895] = '{54.2898453843, 82.2733038412, -77.8072925629, 20.0271688953, 76.7443179736, -33.1412270402, -78.8017580332, -34.978066449};
test_label[361] = '{20.0271688953};
test_output[361] = '{62.2500970993};
############ END DEBUG ############*/
test_input[2896:2903] = '{32'h42a5d41f, 32'hc251fc34, 32'hc1ec0aba, 32'hc2742f21, 32'hc2a61a8f, 32'hc28041ef, 32'hc24bd159, 32'hc21be0be};
test_label[362] = '{32'hc2a61a8f};
test_output[362] = '{32'h4325f757};
/*############ DEBUG ############
test_input[2896:2903] = '{82.9143018584, -52.4962933525, -29.5052367915, -61.0460252241, -83.0518715553, -64.1287746523, -50.9544412342, -38.9694755602};
test_label[362] = '{-83.0518715553};
test_output[362] = '{165.966173414};
############ END DEBUG ############*/
test_input[2904:2911] = '{32'hc28e84fa, 32'h423d8be5, 32'hc2a6723c, 32'h42a1d602, 32'hc1d866dd, 32'h41af2429, 32'h417d7b5f, 32'h42997236};
test_label[363] = '{32'h417d7b5f};
test_output[363] = '{32'h42822e3f};
/*############ DEBUG ############
test_input[2904:2911] = '{-71.2597170918, 47.3866152105, -83.223114226, 80.9179849058, -27.050225639, 21.892656882, 15.8426197811, 76.7230679512};
test_label[363] = '{15.8426197811};
test_output[363] = '{65.0903246648};
############ END DEBUG ############*/
test_input[2912:2919] = '{32'h41e8de99, 32'hc28d0f33, 32'h4287cf22, 32'h42804688, 32'hc2ae6cef, 32'h425807c4, 32'h42b934dc, 32'hc18bd757};
test_label[364] = '{32'hc28d0f33};
test_output[364] = '{32'h43232208};
/*############ DEBUG ############
test_input[2912:2919] = '{29.1086895639, -70.5296873686, 67.9045526964, 64.1377557512, -87.2127574052, 54.0075852677, 92.6032439789, -17.4801467865};
test_label[364] = '{-70.5296873686};
test_output[364] = '{163.132931347};
############ END DEBUG ############*/
test_input[2920:2927] = '{32'h429c43de, 32'hc1fe67ac, 32'hc2345e2c, 32'hc2891820, 32'hc29dd963, 32'hc229da01, 32'h42988a74, 32'hc275eea9};
test_label[365] = '{32'h429c43de};
test_output[365] = '{32'h3e13dc54};
/*############ DEBUG ############
test_input[2920:2927] = '{78.1325514526, -31.8006211883, -45.0919646977, -68.5471221664, -78.9245810751, -42.4628934477, 76.2704161024, -61.483065737};
test_label[365] = '{78.1325514526};
test_output[365] = '{0.144395165833};
############ END DEBUG ############*/
test_input[2928:2935] = '{32'h42a80909, 32'h42b57c8d, 32'hc2b7a095, 32'hc115e4d4, 32'h4277b5f4, 32'hc2998128, 32'hc14eb0fe, 32'h4297ca33};
test_label[366] = '{32'hc2998128};
test_output[366] = '{32'h43277f29};
/*############ DEBUG ############
test_input[2928:2935] = '{84.0176450127, 90.7432595434, -91.813638449, -9.36836618488, 61.9276878138, -76.7522610704, -12.9182108762, 75.8949229864};
test_label[366] = '{-76.7522610704};
test_output[366] = '{167.496720033};
############ END DEBUG ############*/
test_input[2936:2943] = '{32'h42b3645b, 32'hc1147eaa, 32'hc24496da, 32'hc29bed54, 32'hc2230609, 32'h4261757b, 32'hc2a68b1a, 32'hc2405519};
test_label[367] = '{32'hc29bed54};
test_output[367] = '{32'h4327a8d8};
/*############ DEBUG ############
test_input[2936:2943] = '{89.6960068698, -9.28092340036, -49.1473150976, -77.9635349948, -40.7558935883, 56.364727191, -83.2716847695, -48.0831038938};
test_label[367] = '{-77.9635349948};
test_output[367] = '{167.659541865};
############ END DEBUG ############*/
test_input[2944:2951] = '{32'hc212c143, 32'h42ad236d, 32'h4204aac7, 32'h420caa60, 32'h40abaa19, 32'hc28a9c3b, 32'hc289f93e, 32'h410878a0};
test_label[368] = '{32'h4204aac7};
test_output[368] = '{32'h42559c12};
/*############ DEBUG ############
test_input[2944:2951] = '{-36.688732537, 86.5691890306, 33.1667748461, 35.1663818904, 5.36451394676, -69.3051397331, -68.9868018006, 8.52944957856};
test_label[368] = '{33.1667748461};
test_output[368] = '{53.4024141845};
############ END DEBUG ############*/
test_input[2952:2959] = '{32'hc28ae731, 32'hc206fb33, 32'hc234f83d, 32'h42bd3902, 32'h424f5046, 32'h3fea0210, 32'h42c070ad, 32'hc176aa22};
test_label[369] = '{32'h42c070ad};
test_output[369] = '{32'h3e3ad1c2};
/*############ DEBUG ############
test_input[2952:2959] = '{-69.4515484197, -33.7453104196, -45.2424200224, 94.611345499, 51.8283938213, 1.82818791449, 96.2200682304, -15.4165365832};
test_label[369] = '{96.2200682304};
test_output[369] = '{0.182440789162};
############ END DEBUG ############*/
test_input[2960:2967] = '{32'h42bdcf0d, 32'h420b7b18, 32'hc22000b4, 32'h425fd29d, 32'hc28f628d, 32'hc1bb2595, 32'hc20c645c, 32'hc1892297};
test_label[370] = '{32'hc22000b4};
test_output[370] = '{32'h4306e7b4};
/*############ DEBUG ############
test_input[2960:2967] = '{94.9043976924, 34.8702100189, -40.000688133, 55.9556775075, -71.6924813427, -23.3933511801, -35.0980057434, -17.1418904671};
test_label[370] = '{-40.000688133};
test_output[370] = '{134.905085825};
############ END DEBUG ############*/
test_input[2968:2975] = '{32'hc2beded7, 32'h41f88c0b, 32'hc29c214c, 32'hc157edce, 32'hc11373cf, 32'hc19198f4, 32'hc26eaf26, 32'hc1e7347c};
test_label[371] = '{32'h41f88c0b};
test_output[371] = '{32'h80000000};
/*############ DEBUG ############
test_input[2968:2975] = '{-95.4352332058, 31.0683805666, -78.0650325948, -13.4955579299, -9.2157740493, -18.1996847844, -59.6710423255, -28.9006264752};
test_label[371] = '{31.0683805666};
test_output[371] = '{-0.0};
############ END DEBUG ############*/
test_input[2976:2983] = '{32'h42aa5634, 32'h4229ba7e, 32'hc2ab56aa, 32'h3fea523b, 32'h42c7808c, 32'hc2091821, 32'h42b70752, 32'h42a3c29c};
test_label[372] = '{32'h42c7808c};
test_output[372] = '{32'h398b0892};
/*############ DEBUG ############
test_input[2976:2983] = '{85.1683666649, 42.4321195373, -85.6692663854, 1.83063450528, 99.7510645662, -34.2735651561, 91.5142977814, 81.8800974176};
test_label[372] = '{99.7510645662};
test_output[372] = '{0.000265185304816};
############ END DEBUG ############*/
test_input[2984:2991] = '{32'h42880d0e, 32'hc2bd2880, 32'h4205149f, 32'h41840baa, 32'hc281dc74, 32'h41a32c13, 32'hc0ce91fe, 32'h420f0ba8};
test_label[373] = '{32'h41a32c13};
test_output[373] = '{32'h423e8413};
/*############ DEBUG ############
test_input[2984:2991] = '{68.0254991906, -94.579102263, 33.2701388057, 16.5056945343, -64.9305757677, 20.3965208937, -6.45532127439, 35.7613812412};
test_label[373] = '{20.3965208937};
test_output[373] = '{47.6289782969};
############ END DEBUG ############*/
test_input[2992:2999] = '{32'h4227d64b, 32'hc21f7284, 32'h42acf735, 32'h429dedc2, 32'hc26fc93e, 32'h4247535f, 32'h42bdaf25, 32'h42846e44};
test_label[374] = '{32'hc21f7284};
test_output[374] = '{32'h4306b443};
/*############ DEBUG ############
test_input[2992:2999] = '{41.9592695873, -39.8618303389, 86.4828267946, 78.9643673885, -59.946525147, 49.8314169104, 94.8420810994, 66.2153628897};
test_label[374] = '{-39.8618303389};
test_output[374] = '{134.704145757};
############ END DEBUG ############*/
test_input[3000:3007] = '{32'hc04ce4f0, 32'hc1ffc610, 32'h42bc4a3d, 32'h42c2cac1, 32'h41dc483c, 32'hc2684e35, 32'h4292366a, 32'h42b57e7d};
test_label[375] = '{32'h41dc483c};
test_output[375] = '{32'h428bcccb};
/*############ DEBUG ############
test_input[3000:3007] = '{-3.20147332144, -31.9717108161, 94.144996652, 97.3960045114, 27.5352714709, -58.0763724048, 73.1062743813, 90.7470473207};
test_label[375] = '{27.5352714709};
test_output[375] = '{69.8999831002};
############ END DEBUG ############*/
test_input[3008:3015] = '{32'h424e606e, 32'h41d2a79c, 32'hc2b6114a, 32'h4160d868, 32'h4283b44e, 32'hc0de226b, 32'h429b0b8c, 32'h413a9f74};
test_label[376] = '{32'hc2b6114a};
test_output[376] = '{32'h43288e6c};
/*############ DEBUG ############
test_input[3008:3015] = '{51.5941689849, 26.3318409155, -91.0337657763, 14.0528337146, 65.8521547323, -6.94170119754, 77.5225540619, 11.6639294237};
test_label[376] = '{-91.0337657763};
test_output[376] = '{168.556328381};
############ END DEBUG ############*/
test_input[3016:3023] = '{32'h41c81fc0, 32'h42975908, 32'hc27d49f6, 32'hc1bd4d77, 32'hc11fbdea, 32'hc28ee8db, 32'hc29ebaf7, 32'h42c6b72e};
test_label[377] = '{32'hc29ebaf7};
test_output[377] = '{32'h4332b912};
/*############ DEBUG ############
test_input[3016:3023] = '{25.0155030473, 75.6738857777, -63.3222275567, -23.6628250593, -9.98386601025, -71.454794207, -79.3651651314, 99.3577727614};
test_label[377] = '{-79.3651651314};
test_output[377] = '{178.722937893};
############ END DEBUG ############*/
test_input[3024:3031] = '{32'h4140f0ed, 32'h413c58de, 32'h4071539f, 32'hc21657fe, 32'h4129aa94, 32'h424b4106, 32'hc2a1f0a3, 32'h4291c0ea};
test_label[378] = '{32'h413c58de};
test_output[378] = '{32'h42746b9d};
/*############ DEBUG ############
test_input[3024:3031] = '{12.0588195238, 11.7716957211, 3.77072874347, -37.5859287921, 10.6041446273, 50.8135006984, -80.9699967506, 72.876786517};
test_label[378] = '{11.7716957211};
test_output[378] = '{61.1050907961};
############ END DEBUG ############*/
test_input[3032:3039] = '{32'h41f80c34, 32'hc0cc4544, 32'hc228acdb, 32'hc28c359a, 32'hc205d117, 32'h426b1faf, 32'hc2944117, 32'h42789469};
test_label[379] = '{32'hc28c359a};
test_output[379] = '{32'h4304489c};
/*############ DEBUG ############
test_input[3032:3039] = '{31.0059592653, -6.38345543204, -42.1688059366, -70.1046888961, -33.4541907736, 58.7809400896, -74.1271261242, 62.1449309868};
test_label[379] = '{-70.1046888961};
test_output[379] = '{132.283631775};
############ END DEBUG ############*/
test_input[3040:3047] = '{32'h41e66d54, 32'hc2a17f01, 32'h428fe9f3, 32'hc2bc3ec0, 32'h423a1379, 32'hc2159b68, 32'h428af29d, 32'h4209f042};
test_label[380] = '{32'h423a1379};
test_output[380] = '{32'h41cc2513};
/*############ DEBUG ############
test_input[3040:3047] = '{28.8033834071, -80.7480560503, 71.9569355436, -94.1225614149, 46.5190162401, -37.4017628871, 69.473852944, 34.4846268368};
test_label[380] = '{46.5190162401};
test_output[380] = '{25.5181024409};
############ END DEBUG ############*/
test_input[3048:3055] = '{32'h4241ad39, 32'hc29711e5, 32'hc1e48fda, 32'h40265a36, 32'h42bc4b41, 32'h420e7bba, 32'hc080d336, 32'hc1113554};
test_label[381] = '{32'h42bc4b41};
test_output[381] = '{32'h80000000};
/*############ DEBUG ############
test_input[3048:3055] = '{48.4191635629, -75.5349507187, -28.5702403811, 2.59925609079, 94.1469839107, 35.6208271795, -4.02578259996, -9.07551920322};
test_label[381] = '{94.1469839107};
test_output[381] = '{-0.0};
############ END DEBUG ############*/
test_input[3056:3063] = '{32'h42180990, 32'h4285727c, 32'h414639a9, 32'hc2aaf497, 32'h41583e4d, 32'h426941b1, 32'hc18c036e, 32'hc291f57a};
test_label[382] = '{32'hc291f57a};
test_output[382] = '{32'h430bb40a};
/*############ DEBUG ############
test_input[3056:3063] = '{38.0093373179, 66.7236050872, 12.3890768853, -85.4777182024, 13.5152105567, 58.3141534405, -17.5016755768, -72.9794497198};
test_label[382] = '{-72.9794497198};
test_output[382] = '{139.703277534};
############ END DEBUG ############*/
test_input[3064:3071] = '{32'h42401959, 32'h42c06fd7, 32'h42b4bba2, 32'hc1e45ca4, 32'h41bf953c, 32'hc2a5a56c, 32'hc15d0567, 32'hc0e7132b};
test_label[383] = '{32'hc15d0567};
test_output[383] = '{32'h42dc11fc};
/*############ DEBUG ############
test_input[3064:3071] = '{48.0247520741, 96.2184393401, 90.3664685888, -28.545235179, 23.9478674576, -82.8230875428, -13.8138189178, -7.22108971846};
test_label[383] = '{-13.8138189178};
test_output[383] = '{110.035128364};
############ END DEBUG ############*/
test_input[3072:3079] = '{32'hc2977e6d, 32'hc2099d9c, 32'h424b1c49, 32'h41c31092, 32'h42b66517, 32'h4234de97, 32'hc2b599b3, 32'h41007a3f};
test_label[384] = '{32'h41007a3f};
test_output[384] = '{32'h42a655d0};
/*############ DEBUG ############
test_input[3072:3079] = '{-75.7469256827, -34.4039151794, 50.777623888, 24.3830917821, 91.1974444103, 45.2173726825, -90.8001915703, 8.02984482071};
test_label[384] = '{8.02984482071};
test_output[384] = '{83.1675995896};
############ END DEBUG ############*/
test_input[3080:3087] = '{32'hc2676d25, 32'hc1c0c4ef, 32'h42bc7506, 32'hc29b5e2a, 32'hc2511a87, 32'h420e3359, 32'h4231d363, 32'hc21d5a99};
test_label[385] = '{32'hc2511a87};
test_output[385] = '{32'h43128125};
/*############ DEBUG ############
test_input[3080:3087] = '{-57.8565879012, -24.0961590711, 94.2285607953, -77.6839154162, -52.2759060323, 35.5501451261, 44.4564338264, -39.3384733354};
test_label[385] = '{-52.2759060323};
test_output[385] = '{146.504466828};
############ END DEBUG ############*/
test_input[3088:3095] = '{32'hc0945b05, 32'hc0977eec, 32'hc23de92a, 32'hc2bb478a, 32'h42bfe4ac, 32'hc208ec6d, 32'h420ec1b7, 32'h40032f4b};
test_label[386] = '{32'h40032f4b};
test_output[386] = '{32'h42bbcb32};
/*############ DEBUG ############
test_input[3088:3095] = '{-4.63611092257, -4.7342432186, -47.4776986379, -93.6397278022, 95.946623973, -34.2308828706, 35.6891743002, 2.04976160689};
test_label[386] = '{2.04976160689};
test_output[386] = '{93.8968623661};
############ END DEBUG ############*/
test_input[3096:3103] = '{32'h42c198bb, 32'hc2c78471, 32'h41a017a0, 32'hc13cbd9f, 32'hc25f3b1c, 32'hc1dd319d, 32'h4254c9eb, 32'h42c79c2f};
test_label[387] = '{32'hc13cbd9f};
test_output[387] = '{32'h42df4c9a};
/*############ DEBUG ############
test_input[3096:3103] = '{96.7983016311, -99.7586776654, 20.0115354683, -11.7962943822, -55.8077226257, -27.6492245761, 53.1971839426, 99.8050461335};
test_label[387] = '{-11.7962943822};
test_output[387] = '{111.649609029};
############ END DEBUG ############*/
test_input[3104:3111] = '{32'hc250a40f, 32'h423ec64c, 32'h427d2e58, 32'h42c6b26a, 32'h3fab3bae, 32'h41f83d9a, 32'h42aae17e, 32'h42a02ff1};
test_label[388] = '{32'h42aae17e};
test_output[388] = '{32'h415e8762};
/*############ DEBUG ############
test_input[3104:3111] = '{-52.1602128465, 47.6936511688, 63.2952579548, 99.3484654745, 1.33775875245, 31.030079616, 85.440414096, 80.0936344061};
test_label[388] = '{85.440414096};
test_output[388] = '{13.9080522944};
############ END DEBUG ############*/
test_input[3112:3119] = '{32'hc1caa8c7, 32'h42237d4c, 32'hc2b57aea, 32'hc259e328, 32'hc2c3518b, 32'h412de1af, 32'h3f8c04dc, 32'hc2940ebb};
test_label[389] = '{32'hc2b57aea};
test_output[389] = '{32'h43039cc8};
/*############ DEBUG ############
test_input[3112:3119] = '{-25.3324107439, 40.8723607108, -90.7400655741, -54.4718313092, -97.6592651659, 10.8675989186, 1.09389833727, -74.0287730458};
test_label[389] = '{-90.7400655741};
test_output[389] = '{131.612426285};
############ END DEBUG ############*/
test_input[3120:3127] = '{32'h424fccc6, 32'hc2ab213f, 32'hc2593c95, 32'hc21193ac, 32'h42475771, 32'hc2c55d95, 32'h4290b371, 32'hc25b739b};
test_label[390] = '{32'hc25b739b};
test_output[390] = '{32'h42fe6d3f};
/*############ DEBUG ############
test_input[3120:3127] = '{51.9499755312, -85.5649354841, -54.309163053, -36.394211024, 49.835392125, -98.6827768313, 72.3504751991, -54.8628943078};
test_label[390] = '{-54.8628943078};
test_output[390] = '{127.213369508};
############ END DEBUG ############*/
test_input[3128:3135] = '{32'h4083f1c2, 32'h42518f44, 32'hc20b467c, 32'h4147c782, 32'hc1379a74, 32'hc14014a3, 32'h400cd44b, 32'hc268ee0f};
test_label[391] = '{32'h42518f44};
test_output[391] = '{32'h80000000};
/*############ DEBUG ############
test_input[3128:3135] = '{4.12326138557, 52.3899086051, -34.818834285, 12.4862081518, -11.475207987, -12.0050383379, 2.20045734896, -58.2324772393};
test_label[391] = '{52.3899086051};
test_output[391] = '{-0.0};
############ END DEBUG ############*/
test_input[3136:3143] = '{32'hc206d361, 32'hc2695ff8, 32'h421a8053, 32'h42a90b0d, 32'hc2926830, 32'hc22b754f, 32'h41fbe273, 32'hc24bf506};
test_label[392] = '{32'h41fbe273};
test_output[392] = '{32'h425424e1};
/*############ DEBUG ############
test_input[3136:3143] = '{-33.7064264645, -58.3437192204, 38.6253173082, 84.5215867154, -73.2034875106, -42.8645583447, 31.4855709289, -50.9892790023};
test_label[392] = '{31.4855709289};
test_output[392] = '{53.0360157865};
############ END DEBUG ############*/
test_input[3144:3151] = '{32'hc2764333, 32'h4121d701, 32'h4032c32c, 32'h42af4653, 32'h4297afbc, 32'hc2aba12d, 32'hc1941104, 32'h420d9ae2};
test_label[393] = '{32'h4032c32c};
test_output[393] = '{32'h42a9b03b};
/*############ DEBUG ############
test_input[3144:3151] = '{-61.5656238887, 10.1149908108, 2.79316235241, 87.6373516033, 75.8432325301, -85.8147997908, -18.5083083386, 35.401251686};
test_label[393] = '{2.79316235241};
test_output[393] = '{84.8441967997};
############ END DEBUG ############*/
test_input[3152:3159] = '{32'hc2427dfe, 32'hc1c8b86a, 32'h42371c83, 32'h41e914b7, 32'hc2480a21, 32'h421dc7e2, 32'hc256797f, 32'h4283a174};
test_label[394] = '{32'h42371c83};
test_output[394] = '{32'h41a04cc8};
/*############ DEBUG ############
test_input[3152:3159] = '{-48.6230380194, -25.0900463977, 45.7778451339, 29.1351147694, -50.0098902604, 39.4451966564, -53.618647631, 65.81533643};
test_label[394] = '{45.7778451339};
test_output[394] = '{20.0374912981};
############ END DEBUG ############*/
test_input[3160:3167] = '{32'h41b9a6d1, 32'hc2b98664, 32'h42be49f3, 32'h4275bce6, 32'hc17f4a70, 32'h42a48e3f, 32'hc297d5af, 32'h4260cc75};
test_label[395] = '{32'hc17f4a70};
test_output[395] = '{32'h42de3341};
/*############ DEBUG ############
test_input[3160:3167] = '{23.2064541654, -92.7624832061, 95.1444314459, 61.434472009, -15.9556730394, 82.2778232656, -75.9173507815, 56.1996660593};
test_label[395] = '{-15.9556730394};
test_output[395] = '{111.100107068};
############ END DEBUG ############*/
test_input[3168:3175] = '{32'h41f44073, 32'h422828a8, 32'hc2ae876b, 32'h409783d9, 32'hc23c3623, 32'hc2424327, 32'hc2c6aaee, 32'h42458e79};
test_label[396] = '{32'h41f44073};
test_output[396] = '{32'h4196ddcf};
/*############ DEBUG ############
test_input[3168:3175] = '{30.531468801, 42.039701497, -87.2644878077, 4.73484488329, -47.052868367, -48.5655769774, -99.3338475463, 49.3891318047};
test_label[396] = '{30.531468801};
test_output[396] = '{18.8583057621};
############ END DEBUG ############*/
test_input[3176:3183] = '{32'h42ab655c, 32'hc2b62a7e, 32'h42ae99c6, 32'h425f32d2, 32'hc28a080b, 32'h421017aa, 32'h40e5a83d, 32'h42b30c95};
test_label[397] = '{32'hc2b62a7e};
test_output[397] = '{32'h4334bacf};
/*############ DEBUG ############
test_input[3176:3183] = '{85.6979670725, -91.0829908644, 87.3003384702, 55.7996291658, -69.0157113806, 36.0231080745, 7.17678671643, 89.5245721063};
test_label[397] = '{-91.0829908644};
test_output[397] = '{180.729721941};
############ END DEBUG ############*/
test_input[3184:3191] = '{32'h424a9618, 32'hc0bb4e24, 32'h4232ada3, 32'h42c3ceed, 32'h4282e19e, 32'hc15b229f, 32'hc28df913, 32'hc159c6d5};
test_label[398] = '{32'hc0bb4e24};
test_output[398] = '{32'h42cf83cf};
/*############ DEBUG ############
test_input[3184:3191] = '{50.6465776118, -5.85328852103, 44.6695661905, 97.904148947, 65.440657554, -13.6959527397, -70.9864720908, -13.6110432989};
test_label[398] = '{-5.85328852103};
test_output[398] = '{103.757437468};
############ END DEBUG ############*/
test_input[3192:3199] = '{32'h4288e07d, 32'h4213aac5, 32'hc29659a2, 32'h423107de, 32'h41d204de, 32'hc28b575d, 32'hc1ea2129, 32'hc294bcdc};
test_label[399] = '{32'h423107de};
test_output[399] = '{32'h41c17236};
/*############ DEBUG ############
test_input[3192:3199] = '{68.4384514908, 36.9167659538, -75.1750635601, 44.2576841094, 26.2523770817, -69.6706304772, -29.2661916772, -74.3688666321};
test_label[399] = '{44.2576841094};
test_output[399] = '{24.1807673814};
############ END DEBUG ############*/
test_input[3200:3207] = '{32'h42c121cb, 32'hc2c59d88, 32'h41481f68, 32'hc2736aad, 32'h40b801a9, 32'h424816b9, 32'h420e612e, 32'h4161d24f};
test_label[400] = '{32'h4161d24f};
test_output[400] = '{32'h42a4e781};
/*############ DEBUG ############
test_input[3200:3207] = '{96.5659997548, -98.8076746904, 12.5076671743, -60.8541746679, 5.75020246356, 50.0221913067, 35.5949031883, 14.1138447697};
test_label[400] = '{14.1138447697};
test_output[400] = '{82.4521549851};
############ END DEBUG ############*/
test_input[3208:3215] = '{32'hc291a473, 32'h423cba68, 32'hc263743e, 32'hc20b98cf, 32'h41d81dc0, 32'hc2c5601b, 32'h42b861f6, 32'h42801b96};
test_label[401] = '{32'h42b861f6};
test_output[401] = '{32'h2b29a800};
/*############ DEBUG ############
test_input[3208:3215] = '{-72.8211925158, 47.1820358406, -56.8635192247, -34.899226632, 27.0145262069, -98.6877065077, 92.1913303159, 64.0538813359};
test_label[401] = '{92.1913303159};
test_output[401] = '{6.02740080069e-13};
############ END DEBUG ############*/
test_input[3216:3223] = '{32'h428a96e0, 32'h42a8ddc4, 32'hc29f58fc, 32'h42c1e8be, 32'h420f0060, 32'h4286601d, 32'h426cf717, 32'h42363db9};
test_label[402] = '{32'h428a96e0};
test_output[402] = '{32'h41dd4778};
/*############ DEBUG ############
test_input[3216:3223] = '{69.2946806236, 84.4331354838, -79.6737985355, 96.9545736816, 35.7503657891, 67.1877221555, 59.2412990011, 45.5602775545};
test_label[402] = '{69.2946806236};
test_output[402] = '{27.6598967056};
############ END DEBUG ############*/
test_input[3224:3231] = '{32'h4223d45a, 32'h4258489e, 32'hc2b7de82, 32'h42458a95, 32'hc29cf8bd, 32'h42c5bd01, 32'hc2667209, 32'h42543c59};
test_label[403] = '{32'h42c5bd01};
test_output[403] = '{32'h80000000};
/*############ DEBUG ############
test_input[3224:3231] = '{40.9573745329, 54.0709165325, -91.9345865491, 49.3853344772, -78.4858139501, 98.869144704, -57.6113620088, 53.0589319718};
test_label[403] = '{98.869144704};
test_output[403] = '{-0.0};
############ END DEBUG ############*/
test_input[3232:3239] = '{32'hc1db2f3f, 32'hc2aae938, 32'hc2af18b9, 32'hc2a66f55, 32'h4223c54b, 32'hc284b07b, 32'hc2c44d81, 32'hc2bd6c2a};
test_label[404] = '{32'hc1db2f3f};
test_output[404] = '{32'h4288ae75};
/*############ DEBUG ############
test_input[3232:3239] = '{-27.3980694931, -85.4555061499, -87.5482897364, -83.2174456172, 40.9426705854, -66.3446902001, -98.1513728227, -94.7112557433};
test_label[404] = '{-27.3980694931};
test_output[404] = '{68.3407400785};
############ END DEBUG ############*/
test_input[3240:3247] = '{32'h42bd5fe3, 32'h4192d104, 32'h424ccdc0, 32'hc2a9226b, 32'hc1a8f497, 32'hc295e78e, 32'hc2792a7b, 32'hc1ac7abb};
test_label[405] = '{32'h4192d104};
test_output[405] = '{32'h4298aba2};
/*############ DEBUG ############
test_input[3240:3247] = '{94.6872762993, 18.3520581132, 51.2009265674, -84.5672234869, -21.1194285538, -74.9522548055, -62.2914863454, -21.5599276039};
test_label[405] = '{18.3520581132};
test_output[405] = '{76.3352181861};
############ END DEBUG ############*/
test_input[3248:3255] = '{32'hc0a34efe, 32'h423595fd, 32'h41ae5822, 32'hc1122157, 32'h42c7b72f, 32'hc26bd5de, 32'h42236c31, 32'h41b8df11};
test_label[406] = '{32'h42c7b72f};
test_output[406] = '{32'h80000000};
/*############ DEBUG ############
test_input[3248:3255] = '{-5.10339278704, 45.3964714661, 21.7930333485, -9.13313996553, 99.8577766496, -58.9588553005, 40.8556551691, 23.1089199984};
test_label[406] = '{99.8577766496};
test_output[406] = '{-0.0};
############ END DEBUG ############*/
test_input[3256:3263] = '{32'h4200cc1f, 32'hc25c46d7, 32'h4216147b, 32'h4269a405, 32'hc1e7fc4c, 32'h42a11253, 32'h428288a7, 32'h42aec9d5};
test_label[407] = '{32'h42aec9d5};
test_output[407] = '{32'h3a89a0ed};
/*############ DEBUG ############
test_input[3256:3263] = '{32.1993369325, -55.0691793082, 37.5199987885, 58.4101755975, -28.9981920791, 80.5357866564, 65.2669017122, 87.3942049894};
test_label[407] = '{87.3942049894};
test_output[407] = '{0.00105002305652};
############ END DEBUG ############*/
test_input[3264:3271] = '{32'h429d10e6, 32'h42952f24, 32'h425412bc, 32'h42bc18cc, 32'hc29cb99c, 32'h4275ce62, 32'h41f86313, 32'h426f804c};
test_label[408] = '{32'h42bc18cc};
test_output[408] = '{32'h3447fb83};
/*############ DEBUG ############
test_input[3264:3271] = '{78.533002073, 74.5920693503, 53.0182943412, 94.0484314398, -78.3625187861, 61.451547447, 31.0483768981, 59.8752895648};
test_label[408] = '{94.0484314398};
test_output[408] = '{1.86248192338e-07};
############ END DEBUG ############*/
test_input[3272:3279] = '{32'h4044c97f, 32'h42934ac3, 32'h42ab64bf, 32'h427b3ecd, 32'h42b31f47, 32'hc233fe51, 32'hc2537dbd, 32'hc2a7bb02};
test_label[409] = '{32'hc2a7bb02};
test_output[409] = '{32'h432d7275};
/*############ DEBUG ############
test_input[3272:3279] = '{3.07479823601, 73.6460194192, 85.696768211, 62.8113283281, 89.5610863023, -44.9983573003, -52.8727905069, -83.8652504121};
test_label[409] = '{-83.8652504121};
test_output[409] = '{173.447097064};
############ END DEBUG ############*/
test_input[3280:3287] = '{32'h4205646c, 32'hc207f851, 32'hc29b2718, 32'h42134efd, 32'h424500ec, 32'hc1a06125, 32'hc28a864f, 32'h424f4a6f};
test_label[410] = '{32'h42134efd};
test_output[410] = '{32'h41711b56};
/*############ DEBUG ############
test_input[3280:3287] = '{33.3480696248, -33.9924967267, -77.5763574073, 36.8271369221, 49.2509009491, -20.0474344981, -69.2623238824, 51.8226892596};
test_label[410] = '{36.8271369221};
test_output[410] = '{15.0691736552};
############ END DEBUG ############*/
test_input[3288:3295] = '{32'hc2072815, 32'hc2ba0d7e, 32'hc09fa9ca, 32'h421945dc, 32'h42a961fe, 32'hc20a9a1e, 32'hc2b1b39b, 32'hc2993514};
test_label[411] = '{32'hc2993514};
test_output[411] = '{32'h43214b89};
/*############ DEBUG ############
test_input[3288:3295] = '{-33.7891436147, -93.0263538229, -4.98947599852, 38.3182226973, 84.6913929142, -34.6505058806, -88.8507905001, -76.6036668654};
test_label[411] = '{-76.6036668654};
test_output[411] = '{161.29505978};
############ END DEBUG ############*/
test_input[3296:3303] = '{32'h411b5d7f, 32'h42116271, 32'hc1e4432e, 32'h4290c1da, 32'hc1ab027d, 32'h42032e4e, 32'hc238c12a, 32'h42407309};
test_label[412] = '{32'h4290c1da};
test_output[412] = '{32'h2dfe7000};
/*############ DEBUG ############
test_input[3296:3303] = '{9.7103261366, 36.3461332262, -28.5328031808, 72.3786197047, -21.3762144259, 32.7952211518, -46.1886359335, 48.1123406443};
test_label[412] = '{72.3786197047};
test_output[412] = '{2.89261947732e-11};
############ END DEBUG ############*/
test_input[3304:3311] = '{32'hc2b85db4, 32'h41836cb4, 32'hc2c74eb7, 32'hc2c1a1c2, 32'hc240a17e, 32'hc21d0c6b, 32'hc22f1a3a, 32'hc194ec22};
test_label[413] = '{32'hc2c74eb7};
test_output[413] = '{32'h42e829e4};
/*############ DEBUG ############
test_input[3304:3311] = '{-92.1830157864, 16.4280769405, -99.6537427473, -96.8159294525, -48.157707938, -39.2621257146, -43.7756104818, -18.6152995763};
test_label[413] = '{-99.6537427473};
test_output[413] = '{116.081819688};
############ END DEBUG ############*/
test_input[3312:3319] = '{32'h418294c8, 32'hc2372dcd, 32'hc2b549f8, 32'h423f60c7, 32'hc10d1b56, 32'hc2808d5b, 32'h4229cd27, 32'hc24429ce};
test_label[414] = '{32'hc10d1b56};
test_output[414] = '{32'h4262ac41};
/*############ DEBUG ############
test_input[3312:3319] = '{16.3226463681, -45.794725745, -90.6444701885, 47.8445089986, -8.81917416431, -64.2760879343, 42.4503457225, -49.0408235477};
test_label[414] = '{-8.81917416431};
test_output[414] = '{56.6682158946};
############ END DEBUG ############*/
test_input[3320:3327] = '{32'hc29aed3a, 32'hc22b3b73, 32'h42813069, 32'h41eb93e4, 32'hc2a193d8, 32'hc2aa732e, 32'hc215d6f8, 32'h420cffe6};
test_label[415] = '{32'h42813069};
test_output[415] = '{32'h2a4b8000};
/*############ DEBUG ############
test_input[3320:3327] = '{-77.4633303254, -42.8080571764, 64.5945474189, 29.4472119499, -80.7887596268, -85.2249617843, -37.45993063, 35.2499017533};
test_label[415] = '{64.5945474189};
test_output[415] = '{1.80744308409e-13};
############ END DEBUG ############*/
test_input[3328:3335] = '{32'hc2ac17f8, 32'h4214ea95, 32'hc23ddc92, 32'hc2a8996f, 32'h426a9676, 32'h418d4e5c, 32'h42aab445, 32'hc2693734};
test_label[416] = '{32'hc2a8996f};
test_output[416] = '{32'h4329a6da};
/*############ DEBUG ############
test_input[3328:3335] = '{-86.0468165908, 37.2290830427, -47.4654009627, -84.299673878, 58.6469355678, 17.6632605233, 85.3520853071, -58.3039080389};
test_label[416] = '{-84.299673878};
test_output[416] = '{169.651759185};
############ END DEBUG ############*/
test_input[3336:3343] = '{32'h42a91b1b, 32'h4272845c, 32'h41272137, 32'h42c239f3, 32'h421d0005, 32'h42c7fa9d, 32'h41fbedad, 32'h425974d6};
test_label[417] = '{32'h4272845c};
test_output[417] = '{32'h421da8fe};
/*############ DEBUG ############
test_input[3336:3343] = '{84.5529387972, 60.6292560828, 10.4456090626, 97.113181763, 39.2500185191, 99.9894756535, 31.4910522518, 54.3640965069};
test_label[417] = '{60.6292560828};
test_output[417] = '{39.4150328813};
############ END DEBUG ############*/
test_input[3344:3351] = '{32'h426cabb0, 32'h4152d453, 32'hc25fc77a, 32'h42b394e4, 32'h41b3c1a9, 32'hc11dda6c, 32'hc292497b, 32'h40c347a0};
test_label[418] = '{32'hc25fc77a};
test_output[418] = '{32'h4311bc51};
/*############ DEBUG ############
test_input[3344:3351] = '{59.1676647317, 13.176836524, -55.9448009066, 89.7908049352, 22.4695610359, -9.86582573543, -73.143514154, 6.10249319564};
test_label[418] = '{-55.9448009066};
test_output[418] = '{145.735605842};
############ END DEBUG ############*/
test_input[3352:3359] = '{32'h42bc27b4, 32'h42683c62, 32'hc171188b, 32'h429c38aa, 32'h42c46a23, 32'hc2ae662c, 32'hc24b499f, 32'hc2b3b1e6};
test_label[419] = '{32'h42683c62};
test_output[419] = '{32'h4220a83c};
/*############ DEBUG ############
test_input[3352:3359] = '{94.0775464284, 58.0589670342, -15.0684920517, 78.1106699025, 98.2072995007, -87.199552925, -50.8218947149, -89.8474591102};
test_label[419] = '{58.0589670342};
test_output[419] = '{40.1642912967};
############ END DEBUG ############*/
test_input[3360:3367] = '{32'hc2ba586c, 32'hc2be0f8c, 32'hbf2cd437, 32'h4242df17, 32'hc19389fd, 32'hc20c52d5, 32'hc2965cf5, 32'h42677ab9};
test_label[420] = '{32'hbf2cd437};
test_output[420] = '{32'h426a2e25};
/*############ DEBUG ############
test_input[3360:3367] = '{-93.1727009622, -95.0303686496, -0.675113162502, 48.7178624225, -18.442376478, -35.0808905392, -75.1815570787, 57.869845448};
test_label[420] = '{-0.675113162502};
test_output[420] = '{58.5450646142};
############ END DEBUG ############*/
test_input[3368:3375] = '{32'hc29eb37a, 32'h428a419d, 32'h41145bdc, 32'hc27c0bf5, 32'hc28d7a96, 32'hc0a649a5, 32'h429a226f, 32'h4273d301};
test_label[421] = '{32'hc28d7a96};
test_output[421] = '{32'h4313ce9a};
/*############ DEBUG ############
test_input[3368:3375] = '{-79.3505434475, 69.1281486299, 9.27242653104, -63.0116758844, -70.7394260699, -5.1964895828, 77.0672508488, 60.9560569371};
test_label[421] = '{-70.7394260699};
test_output[421] = '{147.807033482};
############ END DEBUG ############*/
test_input[3376:3383] = '{32'h427cd4b0, 32'hc29ae9b7, 32'h429d262e, 32'hc19f8924, 32'hc196e31e, 32'hc28d25a3, 32'hc2ba7116, 32'hc20bf9e9};
test_label[422] = '{32'h427cd4b0};
test_output[422] = '{32'h4175dead};
/*############ DEBUG ############
test_input[3376:3383] = '{63.207703522, -77.456470634, 78.574567391, -19.9419633727, -18.8608975853, -70.5735084011, -93.2208676861, -34.9940536795};
test_label[422] = '{63.207703522};
test_output[422] = '{15.366864081};
############ END DEBUG ############*/
test_input[3384:3391] = '{32'hc29c8f6e, 32'h4271baed, 32'hc0a6aa23, 32'h4104f988, 32'h42b0cdb7, 32'h428aa5ca, 32'hc2883946, 32'h40b780b3};
test_label[423] = '{32'hc29c8f6e};
test_output[423] = '{32'h4326ae93};
/*############ DEBUG ############
test_input[3384:3391] = '{-78.2801357263, 60.4325437265, -5.20826864341, 8.31092077628, 88.401788609, 69.3238059512, -68.1118624289, 5.73446027912};
test_label[423] = '{-78.2801357263};
test_output[423] = '{166.68192434};
############ END DEBUG ############*/
test_input[3392:3399] = '{32'h404fc4ed, 32'h41a393ae, 32'hc2c3553e, 32'h422c3aac, 32'h42151176, 32'h42b947a4, 32'h420d1c2a, 32'h41e755b5};
test_label[424] = '{32'h420d1c2a};
test_output[424] = '{32'h4265731d};
/*############ DEBUG ############
test_input[3392:3399] = '{3.24639444144, 20.4471086843, -97.6664890947, 43.0572960565, 37.2670520452, 92.6399205839, 35.2775036637, 28.9168488565};
test_label[424] = '{35.2775036637};
test_output[424] = '{57.3624169202};
############ END DEBUG ############*/
test_input[3400:3407] = '{32'h42c7cca9, 32'hc27ba430, 32'h42a77b0b, 32'hc19eb4e6, 32'hc2c67bc7, 32'h429ac6ca, 32'h42280b39, 32'h42586944};
test_label[425] = '{32'hc19eb4e6};
test_output[425] = '{32'h42ef79e3};
/*############ DEBUG ############
test_input[3400:3407] = '{99.8997300456, -62.9103390241, 83.7403215974, -19.8383291, -99.2417519966, 77.3882592835, 42.0109578701, 54.1027981881};
test_label[425] = '{-19.8383291};
test_output[425] = '{119.738059242};
############ END DEBUG ############*/
test_input[3408:3415] = '{32'hc0b7a37f, 32'hbf7a4098, 32'hc2442ba3, 32'hc291e9d2, 32'h428050d2, 32'hc248d666, 32'hc2481b91, 32'hc1960d64};
test_label[426] = '{32'hc0b7a37f};
test_output[426] = '{32'h428bcb09};
/*############ DEBUG ############
test_input[3408:3415] = '{-5.73870787816, -0.97754814785, -49.0426151055, -72.9566769313, 64.1578484166, -50.2093717507, -50.0269218864, -18.7565376895};
test_label[426] = '{-5.73870787816};
test_output[426] = '{69.8965562948};
############ END DEBUG ############*/
test_input[3416:3423] = '{32'h429a3c6a, 32'hc203f5b0, 32'h425488ed, 32'h42bdb60c, 32'h4291572a, 32'hc216ea44, 32'hc17e7102, 32'hc0ed0b91};
test_label[427] = '{32'h4291572a};
test_output[427] = '{32'h41b17b88};
/*############ DEBUG ############
test_input[3416:3423] = '{77.1179985629, -32.9899287067, 53.1337154051, 94.8555627438, 72.6702438835, -37.728773516, -15.9025900409, -7.40766196635};
test_label[427] = '{72.6702438835};
test_output[427] = '{22.1853188804};
############ END DEBUG ############*/
test_input[3424:3431] = '{32'hc262813c, 32'hc21ae81b, 32'h4192ca21, 32'h429bccc2, 32'h42747daa, 32'h41835a22, 32'hc2adbc6d, 32'h42afc473};
test_label[428] = '{32'h4192ca21};
test_output[428] = '{32'h428b11f1};
/*############ DEBUG ############
test_input[3424:3431] = '{-56.6262057503, -38.7266665877, 18.3486949421, 77.8999179535, 61.1227178551, 16.4190096528, -86.8680157738, 87.8836871691};
test_label[428] = '{18.3486949421};
test_output[428] = '{69.5350383687};
############ END DEBUG ############*/
test_input[3432:3439] = '{32'hbd5fc2af, 32'hc2b7b768, 32'hc2326d2b, 32'hc2bb253d, 32'h3fae3fb7, 32'hc216135d, 32'h42b9b70b, 32'hc22210ec};
test_label[429] = '{32'hc22210ec};
test_output[429] = '{32'h43055fc0};
/*############ DEBUG ############
test_input[3432:3439] = '{-0.0546290230379, -91.8582158439, -44.6066105339, -93.5727273803, 1.36131936769, -37.5189100934, 92.857501986, -40.5165268877};
test_label[429] = '{-40.5165268877};
test_output[429] = '{133.374028874};
############ END DEBUG ############*/
test_input[3440:3447] = '{32'hc0e8e2aa, 32'h4286caa7, 32'h4280aac8, 32'hc1fb9048, 32'hc25f96ec, 32'h425f0040, 32'hc1a58a60, 32'hc17bb310};
test_label[430] = '{32'hc1a58a60};
test_output[430] = '{32'h42b044a9};
/*############ DEBUG ############
test_input[3440:3447] = '{-7.27766912271, 67.395803816, 64.3335581355, -31.4454500274, -55.8973833773, 55.7502443127, -20.6925653283, -15.7312161197};
test_label[430] = '{-20.6925653283};
test_output[430] = '{88.1340987023};
############ END DEBUG ############*/
test_input[3448:3455] = '{32'h42ae77f6, 32'hc241361b, 32'hc2c259c4, 32'hc211f07b, 32'h42a3e365, 32'h42c732c7, 32'hc16ef776, 32'h42a8d108};
test_label[431] = '{32'h42ae77f6};
test_output[431] = '{32'h4145d68d};
/*############ DEBUG ############
test_input[3448:3455] = '{87.2343005263, -48.3028367629, -97.1753225496, -36.4848429454, 81.94413075, 99.5991767511, -14.9354157426, 84.4082645427};
test_label[431] = '{87.2343005263};
test_output[431] = '{12.3648807648};
############ END DEBUG ############*/
test_input[3456:3463] = '{32'h401ed714, 32'h42b121f8, 32'hc181f723, 32'h42aed8a1, 32'hc2543af6, 32'hc1e2e923, 32'hc0f9debc, 32'hc2250ab2};
test_label[432] = '{32'h42b121f8};
test_output[432] = '{32'h3e8dad14};
/*############ DEBUG ############
test_input[3456:3463] = '{2.48187728788, 88.5663430339, -16.245672238, 87.4231056272, -53.0575774467, -28.363836424, -7.80843916932, -41.2604452769};
test_label[432] = '{88.5663430339};
test_output[432] = '{0.276711094568};
############ END DEBUG ############*/
test_input[3464:3471] = '{32'hc15050bb, 32'hc246307c, 32'hc1f7d629, 32'h42ae6b4f, 32'hc188ac13, 32'h42291737, 32'hc26be941, 32'hc2a1f920};
test_label[433] = '{32'h42ae6b4f};
test_output[433] = '{32'h80000000};
/*############ DEBUG ############
test_input[3464:3471] = '{-13.0197091829, -49.5473484822, -30.9795700849, 87.2095852281, -17.0840196973, 42.2726717288, -58.9777883308, -80.9865746987};
test_label[433] = '{87.2095852281};
test_output[433] = '{-0.0};
############ END DEBUG ############*/
test_input[3472:3479] = '{32'hc2c27634, 32'hc234777b, 32'hc29f4644, 32'h42c46eb4, 32'hc279098c, 32'h41c84b4e, 32'h4152f9b1, 32'hc29714fe};
test_label[434] = '{32'hc234777b};
test_output[434] = '{32'h430f5539};
/*############ DEBUG ############
test_input[3472:3479] = '{-97.2308633412, -45.1166816223, -79.6372370398, 98.2162196692, -62.2593241046, 25.0367691057, 13.1859595594, -75.5409983183};
test_label[434] = '{-45.1166816223};
test_output[434] = '{143.332901292};
############ END DEBUG ############*/
test_input[3480:3487] = '{32'h42b71ed9, 32'h4291ebda, 32'hc2177974, 32'h42bedc84, 32'hc1b5e6c6, 32'hc22bf4cc, 32'hc2a7469c, 32'hc29b2935};
test_label[435] = '{32'hc29b2935};
test_output[435] = '{32'h432d0825};
/*############ DEBUG ############
test_input[3480:3487] = '{91.5602475048, 72.9606446403, -37.8686076007, 95.4306975469, -22.7376831111, -42.9890594989, -83.6379097394, -77.5804793713};
test_label[435] = '{-77.5804793713};
test_output[435] = '{173.031811537};
############ END DEBUG ############*/
test_input[3488:3495] = '{32'h40eda758, 32'hc2bfa16d, 32'hc235339a, 32'h419e628c, 32'h42283b57, 32'h40be1221, 32'hc2ac3176, 32'hc27dbbdb};
test_label[436] = '{32'hc2ac3176};
test_output[436] = '{32'h43002790};
/*############ DEBUG ############
test_input[3488:3495] = '{7.42667789715, -95.8152861109, -45.3003921198, 19.7981185064, 42.0579480038, 5.9397132372, -86.0966005525, -63.4334507675};
test_label[436] = '{-86.0966005525};
test_output[436] = '{128.154548557};
############ END DEBUG ############*/
test_input[3496:3503] = '{32'h42be623d, 32'h40e1aae2, 32'h42061d17, 32'hc1baaee6, 32'h42506ea0, 32'h42930915, 32'h4273cad4, 32'hc2470fb0};
test_label[437] = '{32'h4273cad4};
test_output[437] = '{32'h4208f9a5};
/*############ DEBUG ############
test_input[3496:3503] = '{95.1918679511, 7.05210961075, 33.528406236, -23.3353990503, 52.1080308297, 73.517735039, 60.9480758671, -49.7653186829};
test_label[437] = '{60.9480758671};
test_output[437] = '{34.2437920844};
############ END DEBUG ############*/
test_input[3504:3511] = '{32'hc281e4a6, 32'h42aeaec6, 32'hc1918d22, 32'hc24a5cf0, 32'h42bfccac, 32'hc217bf76, 32'h41a529d5, 32'hc1059a51};
test_label[438] = '{32'hc1059a51};
test_output[438] = '{32'h42d0800f};
/*############ DEBUG ############
test_input[3504:3511] = '{-64.9465789199, 87.3413516123, -18.1939133512, -50.5907601299, 95.8997497591, -37.9369740452, 20.6454266517, -8.35017478104};
test_label[438] = '{-8.35017478104};
test_output[438] = '{104.250116448};
############ END DEBUG ############*/
test_input[3512:3519] = '{32'hc1f2503d, 32'hc24a210b, 32'h42c6a041, 32'hc1960a68, 32'hc25a05f7, 32'h42bb705d, 32'hc2baf949, 32'hc24b888e};
test_label[439] = '{32'h42c6a041};
test_output[439] = '{32'h3b737625};
/*############ DEBUG ############
test_input[3512:3519] = '{-30.2891795929, -50.5322696171, 99.312996727, -18.7550807778, -54.5058260415, 93.7194587111, -93.4868851423, -50.8833544801};
test_label[439] = '{99.312996727};
test_output[439] = '{0.00371492772924};
############ END DEBUG ############*/
test_input[3520:3527] = '{32'h42127603, 32'hc2a449b1, 32'hc2977e2f, 32'h42865789, 32'hc1ca2e71, 32'h425c20ce, 32'hc2b2965f, 32'hc28f5b67};
test_label[440] = '{32'hc28f5b67};
test_output[440] = '{32'h430ad978};
/*############ DEBUG ############
test_input[3520:3527] = '{36.6152452796, -82.1439248512, -75.7464544153, 67.1709658322, -25.2726765344, 55.032036134, -89.2936960453, -71.6785205788};
test_label[440] = '{-71.6785205788};
test_output[440] = '{138.849491758};
############ END DEBUG ############*/
test_input[3528:3535] = '{32'h424fc62d, 32'h428a3e0b, 32'h42790f8f, 32'hc1d2050f, 32'hc2816374, 32'hc26b19f0, 32'h400e4dd3, 32'hc224e7e4};
test_label[441] = '{32'hc2816374};
test_output[441] = '{32'h4305d104};
/*############ DEBUG ############
test_input[3528:3535] = '{51.9435292791, 69.1211777947, 62.2651946365, -26.2524695775, -64.6942415972, -58.7753285142, 2.22349997742, -41.226456874};
test_label[441] = '{-64.6942415972};
test_output[441] = '{133.816472008};
############ END DEBUG ############*/
test_input[3536:3543] = '{32'h3fc429d5, 32'hc2a2a364, 32'hc2996d5b, 32'hc229fa5f, 32'h42594029, 32'hc2af9dc3, 32'hc2a88bc1, 32'h4253874c};
test_label[442] = '{32'hc2a88bc1};
test_output[442] = '{32'h430accd1};
/*############ DEBUG ############
test_input[3536:3543] = '{1.53252655399, -81.3191187071, -76.7135817775, -42.4945020475, 54.3126581318, -87.8081251106, -84.2729532804, 52.882127023};
test_label[442] = '{-84.2729532804};
test_output[442] = '{138.800062781};
############ END DEBUG ############*/
test_input[3544:3551] = '{32'hc2a41ac1, 32'h4280ced0, 32'hc2a6d014, 32'h42b35588, 32'h42c346dc, 32'h40b5c85c, 32'h429463d8, 32'h427dde3a};
test_label[443] = '{32'h40b5c85c};
test_output[443] = '{32'h42b7ea83};
/*############ DEBUG ############
test_input[3544:3551] = '{-82.0522563107, 64.4039290365, -83.4064010458, 89.6670570081, 97.6383957398, 5.68070805073, 74.1950075524, 63.4670195681};
test_label[443] = '{5.68070805073};
test_output[443] = '{91.9580328461};
############ END DEBUG ############*/
test_input[3552:3559] = '{32'hc271b2d5, 32'hc28557a1, 32'h41cebce5, 32'h41207942, 32'hc2a4da5b, 32'hc2a03a7c, 32'hc295b3a3, 32'h3fb1cf11};
test_label[444] = '{32'hc271b2d5};
test_output[444] = '{32'h42ac88a4};
/*############ DEBUG ############
test_input[3552:3559] = '{-60.4246417687, -66.6711498429, 25.8422335911, 10.0296041578, -82.4264732869, -80.1142288968, -74.8508554818, 1.38913171762};
test_label[444] = '{-60.4246417687};
test_output[444] = '{86.2668754956};
############ END DEBUG ############*/
test_input[3560:3567] = '{32'h419c18eb, 32'h41df1524, 32'hc28e1b15, 32'h4148a28e, 32'h42b90938, 32'hc24c577b, 32'hc2a38a61, 32'hc2adbe75};
test_label[445] = '{32'h41df1524};
test_output[445] = '{32'h428143ee};
/*############ DEBUG ############
test_input[3560:3567] = '{19.512167009, 27.8853230551, -71.052896312, 12.5396860322, 92.5180015844, -51.0854308428, -81.7702682764, -86.8719835953};
test_label[445] = '{27.8853230551};
test_output[445] = '{64.6326785292};
############ END DEBUG ############*/
test_input[3568:3575] = '{32'hc1b8c483, 32'h41bf2b57, 32'h424995f4, 32'h4181a6d5, 32'hc2228210, 32'h42462d5d, 32'hc1e8fb64, 32'hc2aaa2e8};
test_label[446] = '{32'hc2228210};
test_output[446] = '{32'h42b6c1e2};
/*############ DEBUG ############
test_input[3568:3575] = '{-23.0959537357, 23.896161342, 50.3964402715, 16.206460287, -40.6270137926, 49.5442997442, -29.1227502265, -85.3181743803};
test_label[446] = '{-40.6270137926};
test_output[446] = '{91.3786786688};
############ END DEBUG ############*/
test_input[3576:3583] = '{32'hc1a50779, 32'h42174cdd, 32'h42847d66, 32'h41f1527f, 32'h421d35a1, 32'h429deaaf, 32'h4190a602, 32'hc2b9856e};
test_label[447] = '{32'hc2b9856e};
test_output[447] = '{32'h432bb80f};
/*############ DEBUG ############
test_input[3576:3583] = '{-20.6286485928, 37.8250635919, 66.244917423, 30.1652812863, 39.3023732718, 78.9583691826, 18.0810583912, -92.7606014232};
test_label[447] = '{-92.7606014232};
test_output[447] = '{171.718973616};
############ END DEBUG ############*/
test_input[3584:3591] = '{32'hc29dc480, 32'hc22c4e41, 32'hc12651ed, 32'hc2829d93, 32'hc0468263, 32'h401b8cc9, 32'h421f9327, 32'h4253515b};
test_label[448] = '{32'h421f9327};
test_output[448] = '{32'h414ef8d2};
/*############ DEBUG ############
test_input[3584:3591] = '{-78.8837872054, -43.0764184718, -10.3950017125, -65.3077629074, -3.10170810558, 2.43046786907, 39.8937048669, 52.8294499537};
test_label[448] = '{39.8937048669};
test_output[448] = '{12.9357474971};
############ END DEBUG ############*/
test_input[3592:3599] = '{32'hc18db9c2, 32'h42b30aac, 32'hc1c67c10, 32'hc279fecf, 32'hc14ed22d, 32'hc28db016, 32'h41cf7022, 32'h42ba1983};
test_label[449] = '{32'h41cf7022};
test_output[449] = '{32'h42864c48};
/*############ DEBUG ############
test_input[3592:3599] = '{-17.7157027723, 89.5208407146, -24.8105770585, -62.498835483, -12.9263127922, -70.8439208505, 25.9297526145, 93.0498254572};
test_label[449] = '{25.9297526145};
test_output[449] = '{67.1489854974};
############ END DEBUG ############*/
test_input[3600:3607] = '{32'h423f7209, 32'h428134e1, 32'hc243f215, 32'hbf460e3f, 32'hc2978a66, 32'hc1ef2334, 32'h42be547f, 32'hc0f02823};
test_label[450] = '{32'h428134e1};
test_output[450] = '{32'h41f47e78};
/*############ DEBUG ############
test_input[3600:3607] = '{47.8613636035, 64.603279457, -48.986407806, -0.77365486223, -75.7703110017, -29.8921896587, 95.1650324522, -7.50489932137};
test_label[450] = '{64.603279457};
test_output[450] = '{30.5617529952};
############ END DEBUG ############*/
test_input[3608:3615] = '{32'h41825b34, 32'h41213e82, 32'hc158aa42, 32'h4222bcad, 32'hc1d31edc, 32'h4206ccfa, 32'h426c1de6, 32'hc1e3d255};
test_label[451] = '{32'h41213e82};
test_output[451] = '{32'h4243ce46};
/*############ DEBUG ############
test_input[3608:3615] = '{16.2945321732, 10.0777610129, -13.541567244, 40.6842555584, -26.390068998, 33.7001716348, 59.0291983589, -28.4777020118};
test_label[451] = '{10.0777610129};
test_output[451] = '{48.9514373568};
############ END DEBUG ############*/
test_input[3616:3623] = '{32'h42ae3685, 32'h4251b9c0, 32'h428a9a19, 32'hc1fedb16, 32'hc23d55b4, 32'hc2814759, 32'h42be9cf3, 32'hc1948c0d};
test_label[452] = '{32'hc23d55b4};
test_output[452] = '{32'h430ea3f8};
/*############ DEBUG ############
test_input[3616:3623] = '{87.1064827617, 52.4313961343, 69.3009698843, -31.8569746266, -47.3336931271, -64.6393523309, 95.3065414568, -18.5683848056};
test_label[452] = '{-47.3336931271};
test_output[452] = '{142.640509184};
############ END DEBUG ############*/
test_input[3624:3631] = '{32'hc28887bd, 32'h3f883205, 32'hc2782305, 32'hc29bd730, 32'hc1c082d5, 32'hc243f610, 32'h4265d74b, 32'h42090dcf};
test_label[453] = '{32'h4265d74b};
test_output[453] = '{32'h2eb95ae0};
/*############ DEBUG ############
test_input[3624:3631] = '{-68.2651159883, 1.06402646145, -62.034199671, -77.9202877998, -24.0638823993, -48.9902968532, 57.4602463739, 34.2634843915};
test_label[453] = '{57.4602463739};
test_output[453] = '{8.42896863453e-11};
############ END DEBUG ############*/
test_input[3632:3639] = '{32'h42af3ef4, 32'h42869a00, 32'h42a192f6, 32'hc2b0d077, 32'h404bb224, 32'h427a79a9, 32'hc20b9d3c, 32'hc17f5815};
test_label[454] = '{32'hc20b9d3c};
test_output[454] = '{32'h42f50e1e};
/*############ DEBUG ############
test_input[3632:3639] = '{87.6229533646, 67.3007830461, 80.7870317418, -88.4071547609, 3.18274785362, 62.6188078099, -34.9035474992, -15.9590040707};
test_label[454] = '{-34.9035474992};
test_output[454] = '{122.527574765};
############ END DEBUG ############*/
test_input[3640:3647] = '{32'hc190dd4f, 32'h428dae1a, 32'h421e47c0, 32'hc17a8465, 32'hc2520ca2, 32'hc2a105fe, 32'h42a9ca05, 32'hc21dc445};
test_label[455] = '{32'h42a9ca05};
test_output[455] = '{32'h35535d95};
/*############ DEBUG ############
test_input[3640:3647] = '{-18.1080610393, 70.8400392522, 39.5700685485, -15.657322756, -52.5123357146, -80.5117053939, 84.894570762, -39.4416707979};
test_label[455] = '{84.894570762};
test_output[455] = '{7.87398074654e-07};
############ END DEBUG ############*/
test_input[3648:3655] = '{32'hc295b759, 32'h41716856, 32'h429fb73c, 32'h42ac64da, 32'hc2ad6354, 32'h41b02e95, 32'hc25bdd21, 32'hc1b02cda};
test_label[456] = '{32'h42ac64da};
test_output[456] = '{32'h3ae7415d};
/*############ DEBUG ############
test_input[3648:3655] = '{-74.858103563, 15.0879730802, 79.8578799715, 86.1969773524, -86.6939987678, 22.022745217, -54.9659476308, -22.0218996857};
test_label[456] = '{86.1969773524};
test_output[456] = '{0.00176433808839};
############ END DEBUG ############*/
test_input[3656:3663] = '{32'h4281dfb9, 32'h41ff618b, 32'h4149ef79, 32'h4204b4d3, 32'h42625bcd, 32'hc11fa386, 32'hc25f9e25, 32'hc29a3657};
test_label[457] = '{32'hc29a3657};
test_output[457] = '{32'h430e0b17};
/*############ DEBUG ############
test_input[3656:3663] = '{64.9369557907, 31.9226278113, 12.6209654695, 33.1765874727, 56.5896494844, -9.97742309672, -55.9044395604, -77.1061307839};
test_label[457] = '{-77.1061307839};
test_output[457] = '{142.043323581};
############ END DEBUG ############*/
test_input[3664:3671] = '{32'h42bb7e2a, 32'hc2c690c6, 32'h421cc661, 32'hc295bd5b, 32'h4282c5bd, 32'h41b223c2, 32'h418fe04b, 32'hc223ffd3};
test_label[458] = '{32'h418fe04b};
test_output[458] = '{32'h42978617};
/*############ DEBUG ############
test_input[3664:3671] = '{93.7464150494, -99.28275882, 39.1937297762, -74.8698378731, 65.3862105859, 22.2674605828, 17.984518658, -40.9998287993};
test_label[458] = '{17.984518658};
test_output[458] = '{75.7618963914};
############ END DEBUG ############*/
test_input[3672:3679] = '{32'h41d68fb9, 32'hc2057e2c, 32'h420f042c, 32'hc1ddafb9, 32'h429cdf2a, 32'hc11b0175, 32'hc25ef4f9, 32'h4208ec49};
test_label[459] = '{32'hc25ef4f9};
test_output[459] = '{32'h43062cd3};
/*############ DEBUG ############
test_input[3672:3679] = '{26.8201764519, -33.3732163142, 35.7540751371, -27.7108023887, 78.4358654309, -9.68785533457, -55.7392320442, 34.2307485574};
test_label[459] = '{-55.7392320442};
test_output[459] = '{134.175097475};
############ END DEBUG ############*/
test_input[3680:3687] = '{32'hc29b9146, 32'hc250ec51, 32'hc262427a, 32'hc02ed725, 32'h42c6c94d, 32'hc2237ff2, 32'hc2c73568, 32'h42bfbe67};
test_label[460] = '{32'hc2c73568};
test_output[460] = '{32'h434706d0};
/*############ DEBUG ############
test_input[3680:3687] = '{-77.7837337518, -52.2307788113, -56.5649173588, -2.73188145205, 99.3931686322, -40.8749448499, -99.6043089343, 95.8718833815};
test_label[460] = '{-99.6043089343};
test_output[460] = '{199.026610469};
############ END DEBUG ############*/
test_input[3688:3695] = '{32'h3fc6a191, 32'h4281546b, 32'hc16daa85, 32'hc11958de, 32'hc25796e7, 32'h4251c5fc, 32'hc1f8e08a, 32'hc258d461};
test_label[461] = '{32'h4251c5fc};
test_output[461] = '{32'h41438b6a};
/*############ DEBUG ############
test_input[3688:3695] = '{1.55180561112, 64.6648758731, -14.8541302924, -9.58419573482, -53.8973645242, 52.4433441982, -31.1096381401, -54.2074015738};
test_label[461] = '{52.4433441982};
test_output[461] = '{12.2215365982};
############ END DEBUG ############*/
test_input[3696:3703] = '{32'hc2689b46, 32'hc289f32c, 32'h420f3f92, 32'h41e4bf21, 32'h422e8890, 32'hc2992e06, 32'hc1038774, 32'h42bcf5d7};
test_label[462] = '{32'hc2992e06};
test_output[462] = '{32'h432b11ee};
/*############ DEBUG ############
test_input[3696:3703] = '{-58.1516346971, -68.9749471401, 35.8120810504, 28.5933243295, 43.6333632918, -76.5898907429, -8.22057005344, 94.4801529637};
test_label[462] = '{-76.5898907429};
test_output[462] = '{171.070043707};
############ END DEBUG ############*/
test_input[3704:3711] = '{32'hc2781846, 32'h42917fed, 32'h42336699, 32'h42737050, 32'h41506691, 32'h42017d06, 32'hc247c2a3, 32'h429f21f4};
test_label[463] = '{32'h42336699};
test_output[463] = '{32'h420ade6e};
/*############ DEBUG ############
test_input[3704:3711] = '{-62.0237044838, 72.74985432, 44.8501918045, 60.8596787136, 13.0250410676, 32.3720940183, -49.9400738689, 79.5663136185};
test_label[463] = '{44.8501918045};
test_output[463] = '{34.717216815};
############ END DEBUG ############*/
test_input[3712:3719] = '{32'h42bb2a3e, 32'h42507561, 32'hc28502ce, 32'h425cc704, 32'h42bc1a2e, 32'hc1e13ef2, 32'h4284b89a, 32'hc2743d91};
test_label[464] = '{32'h4284b89a};
test_output[464] = '{32'h41e169b6};
/*############ DEBUG ############
test_input[3712:3719] = '{93.5825057939, 52.1146259493, -66.5054796637, 55.1943512143, 94.0511319507, -28.155734127, 66.360553273, -61.0601217675};
test_label[464] = '{66.360553273};
test_output[464] = '{28.1766165151};
############ END DEBUG ############*/
test_input[3720:3727] = '{32'h41ed23f2, 32'hc24f33ea, 32'hc2550f55, 32'hc298ea3d, 32'hc188f3a2, 32'hc2649706, 32'hc11340e0, 32'hc284de39};
test_label[465] = '{32'hc2550f55};
test_output[465] = '{32'h42a5d0a7};
/*############ DEBUG ############
test_input[3720:3727] = '{29.642550867, -51.800695821, -53.2649709846, -76.4574949128, -17.1189621459, -57.1474829522, -9.20333835201, -66.4340311326};
test_label[465] = '{-53.2649709846};
test_output[465] = '{82.9075218515};
############ END DEBUG ############*/
test_input[3728:3735] = '{32'hc2988b63, 32'hc2bbb138, 32'h412f7912, 32'h4246822e, 32'h42026643, 32'h42c3e274, 32'hc20da43c, 32'h4171ff23};
test_label[466] = '{32'h4171ff23};
test_output[466] = '{32'h42a5a290};
/*############ DEBUG ############
test_input[3728:3735] = '{-76.2722395299, -93.8461304394, 10.9670578852, 49.6271269941, 32.5998640296, 97.9422905248, -35.4103838829, 15.124788779};
test_label[466] = '{15.124788779};
test_output[466] = '{82.8175017458};
############ END DEBUG ############*/
test_input[3736:3743] = '{32'hc26a39c2, 32'hc2add466, 32'h42300ecd, 32'hc0ff7798, 32'hc2958ac5, 32'h4200f6db, 32'h4135c821, 32'hc16aee9e};
test_label[467] = '{32'hc0ff7798};
test_output[467] = '{32'h424ffdc2};
/*############ DEBUG ############
test_input[3736:3743] = '{-58.5564045047, -86.9148387106, 44.0144534055, -7.98334886187, -74.7710367177, 32.2410711493, 11.3613593536, -14.6832558254};
test_label[467] = '{-7.98334886187};
test_output[467] = '{51.9978099744};
############ END DEBUG ############*/
test_input[3744:3751] = '{32'h428aeecd, 32'h4275a6f8, 32'hc27f1eb7, 32'hc2947972, 32'hc2aa3edb, 32'hc2c30571, 32'h41452c4d, 32'h426a5dc6};
test_label[468] = '{32'h426a5dc6};
test_output[468] = '{32'h412e00b4};
/*############ DEBUG ############
test_input[3744:3751] = '{69.4664093229, 61.413055546, -63.7799945337, -74.2371955224, -85.1227671376, -97.5106293253, 12.3233153714, 58.5915742083};
test_label[468] = '{58.5915742083};
test_output[468] = '{10.87517202};
############ END DEBUG ############*/
test_input[3752:3759] = '{32'hc202e633, 32'hc1154693, 32'hc2a2e00b, 32'hc2a43cd9, 32'hc2928f11, 32'hc26c9d3a, 32'hc2b49fa5, 32'hc2543dda};
test_label[469] = '{32'hc202e633};
test_output[469] = '{32'h41bb291c};
/*############ DEBUG ############
test_input[3752:3759] = '{-32.724802576, -9.32973002546, -81.4375847128, -82.1188466203, -73.279425569, -59.1535403614, -90.3118053022, -53.0604020764};
test_label[469] = '{-32.724802576};
test_output[469] = '{23.3950725506};
############ END DEBUG ############*/
test_input[3760:3767] = '{32'hc21f2cdf, 32'h41c2bc07, 32'h41d21a0e, 32'hc2281d67, 32'h420e744a, 32'hc28e4c63, 32'h413563f5, 32'hc2c5b391};
test_label[470] = '{32'h41d21a0e};
test_output[470] = '{32'h41159d73};
/*############ DEBUG ############
test_input[3760:3767] = '{-39.7938191698, 24.3418111721, 26.2627213773, -42.0287137955, 35.6135617839, -71.14919229, 11.336903203, -98.8507138684};
test_label[470] = '{26.2627213773};
test_output[470] = '{9.35094002149};
############ END DEBUG ############*/
test_input[3768:3775] = '{32'h40505cb0, 32'hc1c694e7, 32'h41a55940, 32'hc2491428, 32'hc20cd432, 32'hc27b0858, 32'h42b0857e, 32'hc25d441f};
test_label[471] = '{32'hc2491428};
test_output[471] = '{32'h430a87c9};
/*############ DEBUG ############
test_input[3768:3775] = '{3.25565712417, -24.8227055964, 20.6685784303, -50.2696855529, -35.2072236907, -62.7581491326, 88.260727064, -55.3165261676};
test_label[471] = '{-50.2696855529};
test_output[471] = '{138.530412617};
############ END DEBUG ############*/
test_input[3776:3783] = '{32'h428e6bab, 32'hc285a035, 32'hc0db875e, 32'hc18cf96b, 32'h42a9202c, 32'hc26b3eaa, 32'hc2a4f4fe, 32'hc24dfa68};
test_label[472] = '{32'h42a9202c};
test_output[472] = '{32'h35d53dc5};
/*############ DEBUG ############
test_input[3776:3783] = '{71.2102855216, -66.8129062841, -6.86027423141, -17.6217868264, 84.5628342914, -58.8111954871, -82.4785033305, -51.4945368781};
test_label[472] = '{84.5628342914};
test_output[472] = '{1.58877136924e-06};
############ END DEBUG ############*/
test_input[3784:3791] = '{32'h425308fe, 32'hc26c034d, 32'hc2b82baf, 32'hc16c41e8, 32'h42198f2d, 32'h40fbdf56, 32'h42b069e5, 32'h4075a32d};
test_label[473] = '{32'h40fbdf56};
test_output[473] = '{32'h42a0abf0};
/*############ DEBUG ############
test_input[3784:3791] = '{52.7587816382, -59.0032242219, -92.0853216291, -14.7660907961, 38.3898201591, 7.87101287252, 88.2068245778, 3.83808439532};
test_label[473] = '{7.87101287252};
test_output[473] = '{80.3358117052};
############ END DEBUG ############*/
test_input[3792:3799] = '{32'hc25bdeaa, 32'h429aa529, 32'h4043e62c, 32'hc1f073cd, 32'hc2b9e086, 32'h417d2e3f, 32'hc29ae7ec, 32'hc1e4a539};
test_label[474] = '{32'h417d2e3f};
test_output[474] = '{32'h4275fec2};
/*############ DEBUG ############
test_input[3792:3799] = '{-54.9674445603, 77.3225757244, 3.06092362095, -30.0565424685, -92.9385193381, 15.8237906897, -77.4529743587, -28.5806742326};
test_label[474] = '{15.8237906897};
test_output[474] = '{61.4987850346};
############ END DEBUG ############*/
test_input[3800:3807] = '{32'hc1c8f005, 32'hc2a7b1c1, 32'hc2bbbcfd, 32'hc2b3b77e, 32'h41cb7cc9, 32'h40c5b248, 32'hc2bc2037, 32'h40ea77ab};
test_label[475] = '{32'hc2bbbcfd};
test_output[475] = '{32'h42ee9c2f};
/*############ DEBUG ############
test_input[3800:3807] = '{-25.1171969791, -83.8471755473, -93.8691159135, -89.8583832012, 25.4359298869, 6.17801303099, -94.0629186899, 7.32710774437};
test_label[475] = '{-93.8691159135};
test_output[475] = '{119.305045818};
############ END DEBUG ############*/
test_input[3808:3815] = '{32'hc283dd11, 32'h428c406f, 32'hc1e299ee, 32'h428fc9ed, 32'h42c738fa, 32'h42375c84, 32'hc0e2bdcf, 32'h408c01ae};
test_label[476] = '{32'h428fc9ed};
test_output[476] = '{32'h41ddbc32};
/*############ DEBUG ############
test_input[3808:3815] = '{-65.9317674992, 70.1258483413, -28.3251604229, 71.8943891926, 99.6112806424, 45.8403465442, -7.08567005442, 4.37520505817};
test_label[476] = '{71.8943891926};
test_output[476] = '{27.7168914498};
############ END DEBUG ############*/
test_input[3816:3823] = '{32'h426a51de, 32'h429ef567, 32'hc1a92c84, 32'h420ac5c1, 32'h423be48a, 32'h40e7ce7b, 32'hc2a2fb2d, 32'h41275727};
test_label[477] = '{32'h429ef567};
test_output[477] = '{32'h30667fb6};
/*############ DEBUG ############
test_input[3816:3823] = '{58.5799465357, 79.4793024491, -21.1467363717, 34.6931179691, 46.9731830448, 7.24395518174, -81.4905774098, 10.4587777843};
test_label[477] = '{79.4793024491};
test_output[477] = '{8.38550007561e-10};
############ END DEBUG ############*/
test_input[3824:3831] = '{32'hbfdde838, 32'hc1a35d87, 32'h423d0661, 32'hc25b8a5d, 32'hc297b776, 32'h4298bf8f, 32'h416b12fa, 32'h426065a9};
test_label[478] = '{32'hc297b776};
test_output[478] = '{32'h43183b83};
/*############ DEBUG ############
test_input[3824:3831] = '{-1.73364925002, -20.4206668187, 47.2562295802, -54.8851192762, -75.8583234627, 76.3741413417, 14.6921328702, 56.0992764301};
test_label[478] = '{-75.8583234627};
test_output[478] = '{152.232464806};
############ END DEBUG ############*/
test_input[3832:3839] = '{32'hc113e435, 32'hc28a0657, 32'hc0f18a7b, 32'h429565a5, 32'hc1f65908, 32'h41500ca2, 32'h417a01b7, 32'hc2136861};
test_label[479] = '{32'h429565a5};
test_output[479] = '{32'h80000000};
/*############ DEBUG ############
test_input[3832:3839] = '{-9.24321471178, -69.0123856107, -7.54815422081, 74.6985270807, -30.793471418, 13.00308428, 15.6254188063, -36.8519308798};
test_label[479] = '{74.6985270807};
test_output[479] = '{-0.0};
############ END DEBUG ############*/
test_input[3840:3847] = '{32'h40b63ebf, 32'hc1a93780, 32'h429a0cea, 32'hc2167b45, 32'hc0ba97da, 32'hc24d3756, 32'h4180e812, 32'hc22528df};
test_label[480] = '{32'hc2167b45};
test_output[480] = '{32'h42e54a8c};
/*############ DEBUG ############
test_input[3840:3847] = '{5.69515927993, -21.1520995401, 77.0252213379, -37.620380006, -5.83103641331, -51.304039109, 16.1133161266, -41.2899144986};
test_label[480] = '{-37.620380006};
test_output[480] = '{114.645601344};
############ END DEBUG ############*/
test_input[3848:3855] = '{32'h42a8f6b0, 32'hc2ba6737, 32'h4296d88f, 32'h42317d6e, 32'h42b5584f, 32'h42ba5659, 32'h428d6b04, 32'h427fb3e3};
test_label[481] = '{32'hc2ba6737};
test_output[481] = '{32'h433a7318};
/*############ DEBUG ############
test_input[3848:3855] = '{84.4818107036, -93.2015930868, 75.4229624173, 44.3724910278, 90.6724814669, 93.1686512446, 70.7090161862, 63.9256718931};
test_label[481] = '{-93.2015930868};
test_output[481] = '{186.449581083};
############ END DEBUG ############*/
test_input[3856:3863] = '{32'h425c12b0, 32'hc24f2afb, 32'h4227125d, 32'h41ccbdff, 32'hc248cfaa, 32'h42809392, 32'hc21490a1, 32'hc26af2d5};
test_label[482] = '{32'hc21490a1};
test_output[482] = '{32'h42cadbef};
/*############ DEBUG ############
test_input[3856:3863] = '{55.0182484348, -51.7919718583, 41.767932595, 25.5927723471, -50.202795068, 64.2882258625, -37.1412406553, -58.7371412992};
test_label[482] = '{-37.1412406553};
test_output[482] = '{101.429560724};
############ END DEBUG ############*/
test_input[3864:3871] = '{32'h428b91a0, 32'h4236b6c6, 32'hc23e1149, 32'hc2956a22, 32'h415322f5, 32'hc10d3e4a, 32'hc2774070, 32'h413f1226};
test_label[483] = '{32'h415322f5};
test_output[483] = '{32'h42625a82};
/*############ DEBUG ############
test_input[3864:3871] = '{69.7844209961, 45.6784888957, -47.5168807232, -74.7072869623, 13.1960347112, -8.82770685167, -61.8129270738, 11.9419311597};
test_label[483] = '{13.1960347112};
test_output[483] = '{56.5883862849};
############ END DEBUG ############*/
test_input[3872:3879] = '{32'h4231ac14, 32'hc1e8d5eb, 32'hc2651f98, 32'hc225b0b6, 32'hc189f5de, 32'h42ba5f5e, 32'h41a6f658, 32'hc19bcce7};
test_label[484] = '{32'h42ba5f5e};
test_output[484] = '{32'h80000000};
/*############ DEBUG ############
test_input[3872:3879] = '{44.4180443552, -29.1044519039, -57.2808518951, -41.4225686063, -17.2450524478, 93.1862625974, 20.8702848585, -19.4750500433};
test_label[484] = '{93.1862625974};
test_output[484] = '{-0.0};
############ END DEBUG ############*/
test_input[3880:3887] = '{32'hc11b6ecb, 32'hc28ff004, 32'hc17b1426, 32'hc1fa24b1, 32'h42c3777d, 32'h421b264a, 32'h418c016a, 32'h40b64335};
test_label[485] = '{32'hc17b1426};
test_output[485] = '{32'h42e2da01};
/*############ DEBUG ############
test_input[3880:3887] = '{-9.71454887713, -71.9687771441, -15.6924194138, -31.2679150013, 97.7333723974, 38.7873902171, 17.5006910221, 5.69570402676};
test_label[485] = '{-15.6924194138};
test_output[485] = '{113.425791811};
############ END DEBUG ############*/
test_input[3888:3895] = '{32'h423b426c, 32'hc1cb5f23, 32'h41ae485a, 32'h411257f6, 32'h42970d71, 32'hc233a307, 32'h42231c84, 32'hc194e10d};
test_label[486] = '{32'h42970d71};
test_output[486] = '{32'h2abf9000};
/*############ DEBUG ############
test_input[3888:3895] = '{46.8148651555, -25.4214534446, 21.7853273818, 9.14647482717, 75.5262503738, -44.9092062474, 40.7778453867, -18.6098876718};
test_label[486] = '{75.5262503738};
test_output[486] = '{3.40283357048e-13};
############ END DEBUG ############*/
test_input[3896:3903] = '{32'h41646fbb, 32'h42b66b42, 32'h42c736fe, 32'hc27d93cd, 32'hc24e3192, 32'hc19fe776, 32'h427ed987, 32'h4152a1c5};
test_label[487] = '{32'h4152a1c5};
test_output[487] = '{32'h42ace2e3};
/*############ DEBUG ############
test_input[3896:3903] = '{14.2772776428, 91.2094868814, 99.6074046827, -63.3943354988, -51.5484084248, -19.988017954, 63.7124272527, 13.1644947462};
test_label[487] = '{13.1644947462};
test_output[487] = '{86.4431352471};
############ END DEBUG ############*/
test_input[3904:3911] = '{32'h4174762a, 32'h42b024a3, 32'hc22c0eab, 32'h429364e9, 32'h41f897d9, 32'hc28d4817, 32'h429526e8, 32'h42b032cf};
test_label[488] = '{32'h4174762a};
test_output[488] = '{32'h4292ffe5};
/*############ DEBUG ############
test_input[3904:3911] = '{15.2788483696, 88.0715535046, -43.0143231034, 73.6970914786, 31.0741439915, -70.6408010089, 74.5759891738, 88.0992389128};
test_label[488] = '{15.2788483696};
test_output[488] = '{73.4997917877};
############ END DEBUG ############*/
test_input[3912:3919] = '{32'h41e912f5, 32'hc21843bb, 32'hc13883cf, 32'hc253dea1, 32'h4279665e, 32'hc259f5eb, 32'h429dbeae, 32'hc1b48eed};
test_label[489] = '{32'hc21843bb};
test_output[489] = '{32'h42e9e08b};
/*############ DEBUG ############
test_input[3912:3919] = '{29.1342573134, -38.0661442722, -11.5321798303, -52.9674119405, 62.3499690597, -54.4901528056, 78.8724196705, -22.5697870505};
test_label[489] = '{-38.0661442722};
test_output[489] = '{116.938564009};
############ END DEBUG ############*/
test_input[3920:3927] = '{32'h42bc000f, 32'hbf9d8a22, 32'hc036f8f5, 32'h4223fad3, 32'hc25d4d55, 32'h42783dfc, 32'h42a18b7d, 32'hc29b6867};
test_label[490] = '{32'hc25d4d55};
test_output[490] = '{32'h4315535d};
/*############ DEBUG ############
test_input[3920:3927] = '{94.0001118416, -1.23077797361, -2.85894505561, 40.9949446901, -55.325518136, 62.0605298603, 80.7724377631, -77.7039104419};
test_label[490] = '{-55.325518136};
test_output[490] = '{149.325631778};
############ END DEBUG ############*/
test_input[3928:3935] = '{32'h41d50635, 32'h42b316dd, 32'hc01a1b30, 32'h4121fe70, 32'hc2c41a5c, 32'hbf54dfbf, 32'h42be88a9, 32'h42c01490};
test_label[491] = '{32'hc01a1b30};
test_output[491] = '{32'h42c5a83b};
/*############ DEBUG ############
test_input[3928:3935] = '{26.6280311795, 89.5446574548, -2.40790939014, 10.1246182811, -98.0514812266, -0.831539075368, 95.2669181527, 96.0401584144};
test_label[491] = '{-2.40790939014};
test_output[491] = '{98.8285743094};
############ END DEBUG ############*/
test_input[3936:3943] = '{32'h416e9ae0, 32'h422ad044, 32'h426fae16, 32'h41981d69, 32'hc28b7624, 32'hc299de15, 32'hc2c26274, 32'h42a22517};
test_label[492] = '{32'h42a22517};
test_output[492] = '{32'h3032f578};
/*############ DEBUG ############
test_input[3936:3943] = '{14.912811546, 42.7033839325, 59.9200046981, 19.0143598152, -69.7307445267, -76.9337566931, -97.1922887903, 81.0724417482};
test_label[492] = '{81.0724417482};
test_output[492] = '{6.51048548618e-10};
############ END DEBUG ############*/
test_input[3944:3951] = '{32'hc2ae0df7, 32'hc253cb6f, 32'h42aa201f, 32'hc0a9783c, 32'h417a47a8, 32'hc1e01f00, 32'h42b6a732, 32'h42bc00c8};
test_label[493] = '{32'hc0a9783c};
test_output[493] = '{32'h42c6ba7a};
/*############ DEBUG ############
test_input[3944:3951] = '{-87.0272762525, -52.9486667209, 85.0627389192, -5.2959268442, 15.6424940263, -28.0151372383, 91.3265556989, 94.0015262888};
test_label[493] = '{-5.2959268442};
test_output[493] = '{99.364214234};
############ END DEBUG ############*/
test_input[3952:3959] = '{32'hc1f38b2d, 32'h42b2389a, 32'h4190ab3c, 32'h429ed99d, 32'hc0d9abb3, 32'h42bc4ab6, 32'hc25b2b7b, 32'hc04fe4aa};
test_label[494] = '{32'h42bc4ab6};
test_output[494] = '{32'h3bd4703d};
/*############ DEBUG ############
test_input[3952:3959] = '{-30.4429578074, 89.1105481624, 18.0836100686, 79.4250280162, -6.80220946124, 94.1459225322, -54.7924620474, -3.24833163031};
test_label[494] = '{94.1459225322};
test_output[494] = '{0.00648310641221};
############ END DEBUG ############*/
test_input[3960:3967] = '{32'hc26dfe8c, 32'h421f2e6c, 32'hc203935e, 32'hc157ef3c, 32'hc27d067f, 32'hc036d4df, 32'hc0296c60, 32'hc2927c7a};
test_label[495] = '{32'h421f2e6c};
test_output[495] = '{32'h80000000};
/*############ DEBUG ############
test_input[3960:3967] = '{-59.4985801894, 39.7953341236, -32.8939124919, -13.4959070395, -63.2563439494, -2.85674258827, -2.647239719, -73.2431175915};
test_label[495] = '{39.7953341236};
test_output[495] = '{-0.0};
############ END DEBUG ############*/
test_input[3968:3975] = '{32'hc292b7d8, 32'h41b8708d, 32'h42c1ba08, 32'hc1baba5c, 32'hc13b72f3, 32'hc0abdb66, 32'h410df2e2, 32'hc25b657f};
test_label[496] = '{32'h410df2e2};
test_output[496] = '{32'h42affbab};
/*############ DEBUG ############
test_input[3968:3975] = '{-73.3590728197, 23.0549559069, 96.8633400467, -23.3409948356, -11.7155633873, -5.37053211778, 8.87179751339, -54.8491182421};
test_label[496] = '{8.87179751339};
test_output[496] = '{87.9915425333};
############ END DEBUG ############*/
test_input[3976:3983] = '{32'hc28f45c3, 32'h40bbf08b, 32'hc2b30f7e, 32'hc191486c, 32'hc1cf5d81, 32'h423f9615, 32'h411ea32a, 32'h41fe247a};
test_label[497] = '{32'hc1cf5d81};
test_output[497] = '{32'h4293a26b};
/*############ DEBUG ############
test_input[3976:3983] = '{-71.6362563022, 5.87311307294, -89.5302611687, -18.160361409, -25.920656436, 47.8965631436, 9.91483458295, 31.7678110194};
test_label[497] = '{-25.920656436};
test_output[497] = '{73.8172196785};
############ END DEBUG ############*/
test_input[3984:3991] = '{32'h4283cd74, 32'h42962ca9, 32'h422712c5, 32'hc2af8f11, 32'hc2b24959, 32'h41b15a14, 32'hc1813cc1, 32'h4299c91d};
test_label[498] = '{32'h422712c5};
test_output[498] = '{32'h420d1b51};
/*############ DEBUG ############
test_input[3984:3991] = '{65.9012757125, 75.0872300653, 41.7683294011, -87.7794278623, -89.1432555806, 22.1689841351, -16.154664069, 76.8928014682};
test_label[498] = '{41.7683294011};
test_output[498] = '{35.2766757207};
############ END DEBUG ############*/
test_input[3992:3999] = '{32'hc28915ed, 32'h42c0ea05, 32'hc252c70e, 32'hc2c2ede3, 32'h429e339f, 32'hc160fe19, 32'hc2a18159, 32'hc26051f5};
test_label[499] = '{32'hc2a18159};
test_output[499] = '{32'h433135af};
/*############ DEBUG ############
test_input[3992:3999] = '{-68.5428235913, 96.457065606, -52.6943878286, -97.4646236898, 79.1008221717, -14.0620358945, -80.7526337028, -56.0800354405};
test_label[499] = '{-80.7526337028};
test_output[499] = '{177.209699338};
############ END DEBUG ############*/
test_input[4000:4007] = '{32'h42848e7f, 32'h425ca389, 32'h42368111, 32'h41bbcd0a, 32'hc19b97c5, 32'hc031624a, 32'hc20b2e45, 32'h421eb977};
test_label[500] = '{32'h42848e7f};
test_output[500] = '{32'h3778e296};
/*############ DEBUG ############
test_input[4000:4007] = '{66.278309587, 55.1597034748, 45.6260396428, 23.4751163219, -19.4491058476, -2.77162404385, -34.7951848829, 39.6811190624};
test_label[500] = '{66.278309587};
test_output[500] = '{1.48347082804e-05};
############ END DEBUG ############*/
test_input[4008:4015] = '{32'hc2a454b2, 32'hc185bb05, 32'hc1bdcba9, 32'h4285ffe6, 32'hc18ddddb, 32'h41e14301, 32'h42468a4d, 32'hc26b5c84};
test_label[501] = '{32'hc18ddddb};
test_output[501] = '{32'h42a9775d};
/*############ DEBUG ############
test_input[4008:4015] = '{-82.1654213393, -16.716318508, -23.724442701, 66.9998035295, -17.7333273202, 28.1577174282, 49.6350584968, -58.8403486761};
test_label[501] = '{-17.7333273202};
test_output[501] = '{84.7331308784};
############ END DEBUG ############*/
test_input[4016:4023] = '{32'hc2303aae, 32'h42b55b50, 32'hbfc1fdd5, 32'h418ef1e3, 32'hc1189f6c, 32'h42168728, 32'hc0014882, 32'h405d43e5};
test_label[502] = '{32'h42b55b50};
test_output[502] = '{32'h80000000};
/*############ DEBUG ############
test_input[4016:4023] = '{-44.0573029227, 90.6783461481, -1.51555878133, 17.8681085888, -9.53892117023, 37.6319875079, -2.02005059641, 3.45726896126};
test_label[502] = '{90.6783461481};
test_output[502] = '{-0.0};
############ END DEBUG ############*/
test_input[4024:4031] = '{32'h42862b85, 32'hc235a52d, 32'h4202fea8, 32'h4260fda0, 32'hc2a7a717, 32'hc2c51403, 32'h42b378c8, 32'h41ae4821};
test_label[503] = '{32'h4202fea8};
test_output[503] = '{32'h4263f2e8};
/*############ DEBUG ############
test_input[4024:4031] = '{67.0850023216, -45.41130537, 32.7486865443, 56.2476788339, -83.8263506525, -98.5390859625, 89.7359014187, 21.7852183602};
test_label[503] = '{32.7486865443};
test_output[503] = '{56.9872148745};
############ END DEBUG ############*/
test_input[4032:4039] = '{32'hc286bd06, 32'h4218201f, 32'h41a83bb6, 32'hc01b3a5a, 32'h42b6bad5, 32'hc2728ed0, 32'hc200336f, 32'h428407b2};
test_label[504] = '{32'h42b6bad5};
test_output[504] = '{32'h2d2c3000};
/*############ DEBUG ############
test_input[4032:4039] = '{-67.3691844992, 38.0313671757, 21.0291555636, -2.4254366083, 91.3649097787, -60.6394635947, -32.0502289919, 66.0150260995};
test_label[504] = '{91.3649097787};
test_output[504] = '{9.78772618514e-12};
############ END DEBUG ############*/
test_input[4040:4047] = '{32'hc1dc1477, 32'hc2a36133, 32'hc2aefd20, 32'h4299e1bc, 32'hc295beb9, 32'hc2915501, 32'hc280617e, 32'h42c1ec6d};
test_label[505] = '{32'h42c1ec6d};
test_output[505] = '{32'h310ab6f5};
/*############ DEBUG ############
test_input[4040:4047] = '{-27.5099930707, -81.6898393341, -87.4943869079, 76.9408901216, -74.8725063666, -72.6660263355, -64.1904158915, 96.9617695557};
test_label[505] = '{96.9617695557};
test_output[505] = '{2.01856409569e-09};
############ END DEBUG ############*/
test_input[4048:4055] = '{32'h41c47bdb, 32'h410e8e71, 32'hc20f7928, 32'h40ae2064, 32'hc215a1eb, 32'h428c5f0b, 32'h3ee8a814, 32'hc1f46a36};
test_label[506] = '{32'h428c5f0b};
test_output[506] = '{32'h80000000};
/*############ DEBUG ############
test_input[4048:4055] = '{24.560475504, 8.90977620539, -35.8683176968, 5.44145383003, -37.4081223504, 70.1856327142, 0.454407327903, -30.5518613977};
test_label[506] = '{70.1856327142};
test_output[506] = '{-0.0};
############ END DEBUG ############*/
test_input[4056:4063] = '{32'h416f44be, 32'h418aa249, 32'hc0a42ab0, 32'hc0e52c2f, 32'hc111c73a, 32'h42c2cadf, 32'h429f8eda, 32'hc2b55449};
test_label[507] = '{32'hc0a42ab0};
test_output[507] = '{32'h42cd0d8a};
/*############ DEBUG ############
test_input[4056:4063] = '{14.9542827707, 17.3292402414, -5.13021087237, -7.16164363394, -9.11113975731, 97.3962306637, 79.7790096546, -90.6646215352};
test_label[507] = '{-5.13021087237};
test_output[507] = '{102.526441558};
############ END DEBUG ############*/
test_input[4064:4071] = '{32'h41905734, 32'h4201d9ca, 32'h41ba02e3, 32'h413b1c21, 32'h42ad1465, 32'h427bf808, 32'h426529b1, 32'h42891109};
test_label[508] = '{32'h4201d9ca};
test_output[508] = '{32'h42584f00};
/*############ DEBUG ############
test_input[4064:4071] = '{18.0425797823, 32.4626827764, 23.2514087575, 11.6943673888, 86.539832546, 62.9922181741, 57.2907143856, 68.533274357};
test_label[508] = '{32.4626827764};
test_output[508] = '{54.0771497848};
############ END DEBUG ############*/
test_input[4072:4079] = '{32'hc2b3be21, 32'h42b6f666, 32'h426408e3, 32'h42a12b7a, 32'hc2318e5b, 32'hbfa87903, 32'h42355108, 32'h429acb28};
test_label[509] = '{32'h42b6f666};
test_output[509] = '{32'h37a1d11c};
/*############ DEBUG ############
test_input[4072:4079] = '{-89.8713432447, 91.481250158, 57.0086784875, 80.5849186803, -44.3890203615, -1.31619297444, 45.3291335744, 77.3967905325};
test_label[509] = '{91.481250158};
test_output[509] = '{1.92900689191e-05};
############ END DEBUG ############*/
test_input[4080:4087] = '{32'h4265c3a6, 32'h421404c6, 32'hc0d7e1b3, 32'h420475b8, 32'hc26698be, 32'h42bc6842, 32'h420ee4f5, 32'hc0b69b4e};
test_label[510] = '{32'h420ee4f5};
test_output[510] = '{32'h4269eb90};
/*############ DEBUG ############
test_input[4080:4087] = '{57.4410642957, 37.0046624496, -6.74630109594, 33.1149578425, -57.6491638219, 94.2036303191, 35.7235904737, -5.70645807859};
test_label[510] = '{35.7235904737};
test_output[510] = '{58.4800398455};
############ END DEBUG ############*/
test_input[4088:4095] = '{32'h408e944c, 32'hc2b48d15, 32'h41fc0728, 32'h427df6bc, 32'hc1b41c4c, 32'h40ab3948, 32'h427abb78, 32'hc23c5891};
test_label[511] = '{32'h427abb78};
test_output[511] = '{32'h3f9698f1};
/*############ DEBUG ############
test_input[4088:4095] = '{4.45560250584, -90.2755523314, 31.5034937837, 63.4909529086, -22.513816584, 5.35074211196, 62.683075727, -47.0864920622};
test_label[511] = '{62.683075727};
test_output[511] = '{1.17654235019};
############ END DEBUG ############*/
test_input[4096:4103] = '{32'hc1b0ed5e, 32'h421739ac, 32'h425a73e5, 32'hc2386f8a, 32'h408175a2, 32'h418e2580, 32'h40a4ce17, 32'h416c4f67};
test_label[512] = '{32'h408175a2};
test_output[512] = '{32'h424a4531};
/*############ DEBUG ############
test_input[4096:4103] = '{-22.1159013638, 37.8063220707, 54.6131780317, -46.1089249309, 4.04560950914, 17.7683107076, 5.15015754808, 14.7693848917};
test_label[512] = '{4.04560950914};
test_output[512] = '{50.5675685728};
############ END DEBUG ############*/
test_input[4104:4111] = '{32'hc2a2e5f8, 32'hc14a4cd5, 32'hc2633f8a, 32'h41df4e21, 32'h4263868c, 32'hc2080669, 32'hc2a4347d, 32'hc2c1b2e4};
test_label[513] = '{32'hc2a2e5f8};
test_output[513] = '{32'h430a549f};
/*############ DEBUG ############
test_input[4104:4111] = '{-81.4491563788, -12.643757514, -56.8120485476, 27.9131489625, 56.8813929404, -34.0062600999, -82.1025177453, -96.8493948358};
test_label[513] = '{-81.4491563788};
test_output[513] = '{138.330549319};
############ END DEBUG ############*/
test_input[4112:4119] = '{32'hc23c71c4, 32'h42b3ca87, 32'hbfe5438e, 32'hc12daff7, 32'h41ff2cba, 32'hc0c61515, 32'hc2c26409, 32'h42667602};
test_label[514] = '{32'hc0c61515};
test_output[514] = '{32'h42c02bd8};
/*############ DEBUG ############
test_input[4112:4119] = '{-47.1110975328, 89.8955587911, -1.79112411538, -10.8554600454, 31.8968385659, -6.190073531, -97.1953846645, 57.6152414177};
test_label[514] = '{-6.190073531};
test_output[514] = '{96.0856323221};
############ END DEBUG ############*/
test_input[4120:4127] = '{32'hc19d9f75, 32'hc2aa65f6, 32'h4219c661, 32'hc08cea1d, 32'hc250a358, 32'h3fb24b69, 32'h3fcec349, 32'hc266c52f};
test_label[515] = '{32'h3fcec349};
test_output[515] = '{32'h42135047};
/*############ DEBUG ############
test_input[4120:4127] = '{-19.7028599695, -85.1991386887, 38.4437288901, -4.40357808035, -52.1595159613, 1.39292631523, 1.61533462445, -57.6925603807};
test_label[515] = '{1.61533462445};
test_output[515] = '{36.8283942656};
############ END DEBUG ############*/
test_input[4128:4135] = '{32'hc27f835e, 32'h41d3bf8d, 32'h406b0452, 32'h42942a4e, 32'hc2a912dc, 32'h42ad276f, 32'h4175b801, 32'h4219e805};
test_label[516] = '{32'h406b0452};
test_output[516] = '{32'h42a5cf4d};
/*############ DEBUG ############
test_input[4128:4135] = '{-63.8782898094, 26.4685309565, 3.67213862693, 74.0826257757, -84.5368363699, 86.5770191274, 15.3574227935, 38.4765819517};
test_label[516] = '{3.67213862693};
test_output[516] = '{82.904884248};
############ END DEBUG ############*/
test_input[4136:4143] = '{32'hc29276c2, 32'hc2bf373b, 32'h42037277, 32'h42a5f5de, 32'hc1fa9c06, 32'hc232eaa2, 32'hc2541dff, 32'h42a3a0c1};
test_label[517] = '{32'hc2bf373b};
test_output[517] = '{32'h4332dbfa};
/*############ DEBUG ############
test_input[4136:4143] = '{-73.2319460046, -95.6078696245, 32.8617833197, 82.9802089898, -31.3261823773, -44.7291350875, -53.0292939913, 81.8139711061};
test_label[517] = '{-95.6078696245};
test_output[517] = '{178.859278176};
############ END DEBUG ############*/
test_input[4144:4151] = '{32'h41197c37, 32'hc1e17845, 32'h42aed9f1, 32'hc1251fd5, 32'h42908d90, 32'hc288aaf3, 32'h426e6e0c, 32'h42866ef6};
test_label[518] = '{32'h41197c37};
test_output[518] = '{32'h429baa6a};
/*############ DEBUG ############
test_input[4144:4151] = '{9.59282631, -28.1837249795, 87.4256651991, -10.3202716164, 72.2764882133, -68.3338864418, 59.6074693364, 67.2167206657};
test_label[518] = '{9.59282631};
test_output[518] = '{77.8328391543};
############ END DEBUG ############*/
test_input[4152:4159] = '{32'hc28bf8ae, 32'h421b597c, 32'h3f807197, 32'hc23cb5a6, 32'h42282692, 32'hc22de3f1, 32'h42b9a462, 32'hc241f456};
test_label[519] = '{32'h421b597c};
test_output[519] = '{32'h4257ef48};
/*############ DEBUG ############
test_input[4152:4159] = '{-69.9857058238, 38.8373881695, 1.00346650503, -47.1773917157, 42.0376679868, -43.4726001616, 92.8210627131, -48.4886111822};
test_label[519] = '{38.8373881695};
test_output[519] = '{53.9836745436};
############ END DEBUG ############*/
test_input[4160:4167] = '{32'hc2c374eb, 32'h42c52b9c, 32'h41a738d5, 32'hc2a7a683, 32'h42597a40, 32'hc2bb842b, 32'hc169e931, 32'h42341c4b};
test_label[520] = '{32'hc2c374eb};
test_output[520] = '{32'h43445044};
/*############ DEBUG ############
test_input[4160:4167] = '{-97.7283577042, 98.5851767499, 20.9027497152, -83.8252192688, 54.3693859379, -93.7581406095, -14.6194314901, 45.0276315564};
test_label[520] = '{-97.7283577042};
test_output[520] = '{196.313534454};
############ END DEBUG ############*/
test_input[4168:4175] = '{32'hc227f732, 32'hc2b6036b, 32'h41201ee7, 32'h4295ba19, 32'hc2b7fc0e, 32'h419aaf5c, 32'h3f4e7aea, 32'hc1c6319b};
test_label[521] = '{32'hc2b6036b};
test_output[521] = '{32'h4325dec2};
/*############ DEBUG ############
test_input[4168:4175] = '{-41.9914015954, -91.0066775565, 10.0075441218, 74.8634732931, -91.9922907388, 19.3356242196, 0.806563000087, -24.7742215927};
test_label[521] = '{-91.0066775565};
test_output[521] = '{165.87015085};
############ END DEBUG ############*/
test_input[4176:4183] = '{32'hc152785f, 32'h42bcb376, 32'h42ad4972, 32'hc1537b1f, 32'hc1255e7e, 32'h4210df04, 32'hc28cc584, 32'h427576d9};
test_label[522] = '{32'hc152785f};
test_output[522] = '{32'h42d702bd};
/*############ DEBUG ############
test_input[4176:4183] = '{-13.154387624, 94.350509966, 86.6434440784, -13.2175589045, -10.3355698279, 36.2177878522, -70.3857740413, 61.3660614199};
test_label[522] = '{-13.154387624};
test_output[522] = '{107.505347128};
############ END DEBUG ############*/
test_input[4184:4191] = '{32'h40eee5ac, 32'hc19740fe, 32'hc2863622, 32'h42782664, 32'hc1802b94, 32'hc2c747aa, 32'hc2a55eff, 32'hc249bbc2};
test_label[523] = '{32'hc2a55eff};
test_output[523] = '{32'h4310b919};
/*############ DEBUG ############
test_input[4184:4191] = '{7.46553618409, -18.9067340822, -67.1057299743, 62.0374895433, -16.0212788389, -99.6399685531, -82.6855418808, -50.433358317};
test_label[523] = '{-82.6855418808};
test_output[523] = '{144.723031424};
############ END DEBUG ############*/
test_input[4192:4199] = '{32'h3f91af79, 32'hc27d469d, 32'hc24e7c0b, 32'hc23a76bf, 32'hc19569cb, 32'hc2319f4a, 32'hc2b42301, 32'hc26be1ee};
test_label[524] = '{32'h3f91af79};
test_output[524] = '{32'h312a749d};
/*############ DEBUG ############
test_input[4192:4199] = '{1.1381674925, -63.3189588192, -51.6211352108, -46.6159624883, -18.6766567015, -44.4055542537, -90.068365314, -58.9706341187};
test_label[524] = '{1.1381674925};
test_output[524] = '{2.48045417847e-09};
############ END DEBUG ############*/
test_input[4200:4207] = '{32'h4259a129, 32'hc29fc828, 32'hc274b203, 32'h424eb5de, 32'h42c529ca, 32'h428aafdb, 32'hc2a3f948, 32'h428adc4b};
test_label[525] = '{32'hc2a3f948};
test_output[525] = '{32'h43349189};
/*############ DEBUG ############
test_input[4200:4207] = '{54.4073847168, -79.890930744, -61.1738377853, 51.6776055362, 98.5816164017, 69.3434698142, -81.9868752724, 69.4302603864};
test_label[525] = '{-81.9868752724};
test_output[525] = '{180.568491674};
############ END DEBUG ############*/
test_input[4208:4215] = '{32'h4204977a, 32'hc2899d03, 32'hc2029f42, 32'hc2c3e4d8, 32'h4266762c, 32'h428b952f, 32'hc25c2194, 32'hc2b73ae9};
test_label[526] = '{32'hc2c3e4d8};
test_output[526] = '{32'h4327bd04};
/*############ DEBUG ############
test_input[4208:4215] = '{33.1479263435, -68.8066631712, -32.6555264598, -97.94695949, 57.615402577, 69.7913739711, -55.0327913778, -91.6150612142};
test_label[526] = '{-97.94695949};
test_output[526] = '{167.738338614};
############ END DEBUG ############*/
test_input[4216:4223] = '{32'hc1c14850, 32'h414e15f7, 32'hc1e2c9d6, 32'hc2b4d680, 32'h42b8e835, 32'h415a7a93, 32'h420f408e, 32'hc038c7db};
test_label[527] = '{32'hc1e2c9d6};
test_output[527] = '{32'h42f19aaa};
/*############ DEBUG ############
test_input[4216:4223] = '{-24.1603092434, 12.8803624587, -28.348552986, -90.4189481247, 92.4535288186, 13.6549253322, 35.8130426754, -2.88719823563};
test_label[527] = '{-28.348552986};
test_output[527] = '{120.802081805};
############ END DEBUG ############*/
test_input[4224:4231] = '{32'h4297bad3, 32'h427d5d87, 32'h42b90ac4, 32'h409ad31a, 32'h426a3458, 32'h4288fe0c, 32'hc296e2a2, 32'h4287bda9};
test_label[528] = '{32'h409ad31a};
test_output[528] = '{32'h42af5d93};
/*############ DEBUG ############
test_input[4224:4231] = '{75.8648944012, 63.3413361845, 92.5210291873, 4.83826929986, 58.5511155267, 68.4961818438, -75.4426430369, 67.8704297268};
test_label[528] = '{4.83826929986};
test_output[528] = '{87.6827599459};
############ END DEBUG ############*/
test_input[4232:4239] = '{32'hc298f6df, 32'hc2c5da1f, 32'hc23a7b85, 32'hc27578e8, 32'hc224935b, 32'hc2c6ad15, 32'h41bd5540, 32'h42b2125f};
test_label[529] = '{32'hc23a7b85};
test_output[529] = '{32'h4307a811};
/*############ DEBUG ############
test_input[4232:4239] = '{-76.4821722418, -98.9260147773, -46.6206249984, -61.3680720818, -41.143901086, -99.3380513855, 23.6666266284, 89.0358844497};
test_label[529] = '{-46.6206249984};
test_output[529] = '{135.656509448};
############ END DEBUG ############*/
test_input[4240:4247] = '{32'h4282967f, 32'hc2a0af0c, 32'hc28ae56d, 32'h41f008aa, 32'hc2222d74, 32'hc193ce74, 32'h3fee0b2e, 32'hc1d2b47b};
test_label[530] = '{32'hc28ae56d};
test_output[530] = '{32'h4306bdf6};
/*############ DEBUG ############
test_input[4240:4247] = '{65.2939365796, -80.3418893598, -69.4481001943, 30.0042295682, -40.5443891602, -18.4758075155, 1.85971616828, -26.3381243676};
test_label[530] = '{-69.4481001943};
test_output[530] = '{134.742036774};
############ END DEBUG ############*/
test_input[4248:4255] = '{32'hc2aea1e8, 32'hc22b0a5f, 32'hc213fb34, 32'h42084a1f, 32'hc2a8ad56, 32'h42b83037, 32'hc2b79650, 32'hc2a6a108};
test_label[531] = '{32'h42084a1f};
test_output[531] = '{32'h4268164f};
/*############ DEBUG ############
test_input[4248:4255] = '{-87.3162215276, -42.7601298914, -36.9953141186, 34.0723824131, -84.3385451441, 92.0941673327, -91.7935796159, -83.3145115202};
test_label[531] = '{34.0723824131};
test_output[531] = '{58.0217849196};
############ END DEBUG ############*/
test_input[4256:4263] = '{32'hc2679f91, 32'h412f61ed, 32'h428fb65a, 32'h4154b6b7, 32'h42bdf996, 32'h429a7a7c, 32'hc19047bd, 32'hc1bb8816};
test_label[532] = '{32'h42bdf996};
test_output[532] = '{32'h32a90ce4};
/*############ DEBUG ############
test_input[4256:4263] = '{-57.9058265693, 10.9614074845, 71.8561541155, 13.2946079457, 94.9874717686, 77.2392282824, -18.0350284934, -23.4414491438};
test_label[532] = '{94.9874717686};
test_output[532] = '{1.96800513379e-08};
############ END DEBUG ############*/
test_input[4264:4271] = '{32'hc156d06b, 32'h428d172c, 32'hbf8bf669, 32'hc26d1b51, 32'hc2b154c7, 32'h40a7432e, 32'hc2b46097, 32'hc19f3dc1};
test_label[533] = '{32'hbf8bf669};
test_output[533] = '{32'h428f4706};
/*############ DEBUG ############
test_input[4264:4271] = '{-13.4258832047, 70.5452573661, -1.09345730753, -59.2766761278, -88.6655814574, 5.2269505037, -90.1886527955, -19.9051542262};
test_label[533] = '{-1.09345730753};
test_output[533] = '{71.6387146736};
############ END DEBUG ############*/
test_input[4272:4279] = '{32'hc223ac6d, 32'hc21710e7, 32'h424d5f43, 32'h42a2f72e, 32'h42585da1, 32'hc2bc4084, 32'h42b17f57, 32'hc1ed8030};
test_label[534] = '{32'hc2bc4084};
test_output[534] = '{32'h4336e01b};
/*############ DEBUG ############
test_input[4272:4279] = '{-40.9183857622, -37.7665051241, 51.3430281613, 81.4827728331, 54.0914326892, -94.1260055196, 88.7487138398, -29.6875913109};
test_label[534] = '{-94.1260055196};
test_output[534] = '{182.875418058};
############ END DEBUG ############*/
test_input[4280:4287] = '{32'hc29d6be5, 32'hc228d2c5, 32'h41576b49, 32'h428a1565, 32'hc25bcace, 32'h41c9b9d5, 32'h4207527b, 32'h41f1aee2};
test_label[535] = '{32'h41f1aee2};
test_output[535] = '{32'h421b5358};
/*############ DEBUG ############
test_input[4280:4287] = '{-78.7107318799, -42.2058304339, 13.4636931368, 69.0417832688, -54.9480508446, 25.2157387001, 33.8305477091, 30.2103913763};
test_label[535] = '{30.2103913763};
test_output[535] = '{38.8313918925};
############ END DEBUG ############*/
test_input[4288:4295] = '{32'h420ddbb2, 32'hc28e85c8, 32'hc29cdef0, 32'h41d91661, 32'h40840c85, 32'h41d63a9c, 32'h4240b98d, 32'h415e16e1};
test_label[536] = '{32'h420ddbb2};
test_output[536] = '{32'h414b7770};
/*############ DEBUG ############
test_input[4288:4295] = '{35.4645446249, -71.2612943308, -78.435424448, 27.1359279067, 4.12652847824, 26.7786177991, 48.1812015236, 13.8805852305};
test_label[536] = '{35.4645446249};
test_output[536] = '{12.7166599006};
############ END DEBUG ############*/
test_input[4296:4303] = '{32'hc2726cfd, 32'hc2a54a07, 32'h41dcd0a8, 32'h4041c0b2, 32'h40a1df0e, 32'h42b02a2b, 32'hc2aa66f1, 32'hc23ec918};
test_label[537] = '{32'h40a1df0e};
test_output[537] = '{32'h42a60c3a};
/*############ DEBUG ############
test_input[4296:4303] = '{-60.6064336682, -82.6445845014, 27.6018837031, 3.02738611827, 5.05847859287, 88.0823613776, -85.2010586741, -47.6963813521};
test_label[537] = '{5.05847859287};
test_output[537] = '{83.0238827847};
############ END DEBUG ############*/
test_input[4304:4311] = '{32'hc294af59, 32'hc2c4acaa, 32'hc257e12c, 32'hc2c0d967, 32'hc281eb4a, 32'h41cd9195, 32'hc2afde42, 32'h42546f7b};
test_label[538] = '{32'hc281eb4a};
test_output[538] = '{32'h42ec2308};
/*############ DEBUG ############
test_input[4304:4311] = '{-74.3424775281, -98.3372324772, -53.9698942568, -96.4246103268, -64.959552701, 25.6960844805, -87.9340970003, 53.1088661344};
test_label[538] = '{-64.959552701};
test_output[538] = '{118.068418835};
############ END DEBUG ############*/
test_input[4312:4319] = '{32'h410069fa, 32'h4282ab7e, 32'h429162f0, 32'hc287f453, 32'h421019ab, 32'h42495967, 32'hc2ad0581, 32'hc2ba3db9};
test_label[539] = '{32'hc2ad0581};
test_output[539] = '{32'h431f3462};
/*############ DEBUG ############
test_input[4312:4319] = '{8.02587275664, 65.3349486448, 72.6932338545, -67.9771991135, 36.0250656281, 50.3373061585, -86.5107498743, -93.1205541777};
test_label[539] = '{-86.5107498743};
test_output[539] = '{159.204620816};
############ END DEBUG ############*/
test_input[4320:4327] = '{32'hc29df42f, 32'hc29eec6b, 32'h4274d1eb, 32'h42c588f6, 32'h42b02ab2, 32'h4227a77d, 32'h41e02ee8, 32'h41e603bb};
test_label[540] = '{32'h42b02ab2};
test_output[540] = '{32'h412af235};
/*############ DEBUG ############
test_input[4320:4327] = '{-78.976924821, -79.4617519333, 61.2049976354, 98.7674992159, 88.0833900144, 41.9135628795, 28.0229035039, 28.7518205833};
test_label[540] = '{88.0833900144};
test_output[540] = '{10.6841321074};
############ END DEBUG ############*/
test_input[4328:4335] = '{32'h40da4e7e, 32'h425d624e, 32'h429ae9a3, 32'h42317202, 32'hc2ab1d4c, 32'hc0ed3e86, 32'hc1a4d9a4, 32'h41a59eae};
test_label[541] = '{32'hc2ab1d4c};
test_output[541] = '{32'h43230378};
/*############ DEBUG ############
test_input[4328:4335] = '{6.82208135376, 55.3460007516, 77.4563220389, 44.361335476, -85.5572221469, -7.4138822621, -20.6062698114, 20.7024797569};
test_label[541] = '{-85.5572221469};
test_output[541] = '{163.013544186};
############ END DEBUG ############*/
test_input[4336:4343] = '{32'h418bcdb1, 32'h419161be, 32'hc1a76871, 32'h3fe831e7, 32'hc2a9ab0f, 32'h42408d58, 32'h42a7c77b, 32'h41fd7f0a};
test_label[542] = '{32'h419161be};
test_output[542] = '{32'h42836f0c};
/*############ DEBUG ############
test_input[4336:4343] = '{17.4754349003, 18.1727255257, -20.9259959714, 1.81402286056, -84.8340952887, 48.1380312028, 83.8896128678, 31.6870312899};
test_label[542] = '{18.1727255257};
test_output[542] = '{65.7168873421};
############ END DEBUG ############*/
test_input[4344:4351] = '{32'hc28c7221, 32'h42357ac4, 32'hc13d1231, 32'h40f1e24c, 32'hc2669165, 32'hc25a6af5, 32'h4216dc65, 32'hc28e86a4};
test_label[543] = '{32'hc28c7221};
test_output[543] = '{32'h42e72fc1};
/*############ DEBUG ############
test_input[4344:4351] = '{-70.2229077786, 45.3698877551, -11.8169417233, 7.55887424916, -57.6419855309, -54.6044514195, 37.7152293082, -71.2629715727};
test_label[543] = '{-70.2229077786};
test_output[543] = '{115.593269253};
############ END DEBUG ############*/
test_input[4352:4359] = '{32'h42c4444a, 32'h42291454, 32'hc11466ab, 32'h41246f57, 32'h426d85b1, 32'h42415b1e, 32'h420ddc11, 32'hc2366b31};
test_label[544] = '{32'hc2366b31};
test_output[544] = '{32'h430fbcf1};
/*############ DEBUG ############
test_input[4352:4359] = '{98.1333787169, 42.2698498086, -9.27506494712, 10.2771822983, 59.3805582735, 48.3389830892, 35.4649083231, -45.6046786403};
test_label[544] = '{-45.6046786403};
test_output[544] = '{143.738057357};
############ END DEBUG ############*/
test_input[4360:4367] = '{32'hc25894e8, 32'h429b4e2c, 32'h42c4a46c, 32'h42046b28, 32'h42c4dc41, 32'h429a91de, 32'h41d7e536, 32'h41bcb336};
test_label[545] = '{32'h429a91de};
test_output[545] = '{32'h41ae487e};
/*############ DEBUG ############
test_input[4360:4367] = '{-54.1454176025, 77.6526774733, 98.3211376774, 33.104646547, 98.4301817718, 77.2848952787, 26.9869188512, 23.5875056254};
test_label[545] = '{77.2848952787};
test_output[545] = '{21.7853972183};
############ END DEBUG ############*/
test_input[4368:4375] = '{32'h421b209f, 32'h3e648461, 32'h41b89d86, 32'h42a01ad5, 32'h40f79e41, 32'h424d195a, 32'h41fe1fed, 32'h41a34d6b};
test_label[546] = '{32'h421b209f};
test_output[546] = '{32'h4225150b};
/*############ DEBUG ############
test_input[4368:4375] = '{38.7818564723, 0.223161241324, 23.0769161442, 80.0524063597, 7.73806810818, 51.2747582403, 31.7655884529, 20.4128017192};
test_label[546] = '{38.7818564723};
test_output[546] = '{41.2705498874};
############ END DEBUG ############*/
test_input[4376:4383] = '{32'h401bc2f2, 32'h42bf6db5, 32'h426e0cd3, 32'h419e2253, 32'hbfd66850, 32'h4263446a, 32'h424b0830, 32'h4118a591};
test_label[547] = '{32'hbfd66850};
test_output[547] = '{32'h42c2c756};
/*############ DEBUG ############
test_input[4376:4383] = '{2.433773532, 95.7142692812, 59.5125232532, 19.7667590943, -1.67505834818, 56.8168121429, 50.7579971459, 9.54042165854};
test_label[547] = '{-1.67505834818};
test_output[547] = '{97.3893276294};
############ END DEBUG ############*/
test_input[4384:4391] = '{32'h41b8a8e9, 32'h41255818, 32'hc19c2e48, 32'h4209db83, 32'h41af2e2c, 32'hc21a2dad, 32'h428e73ce, 32'hc2afc19f};
test_label[548] = '{32'h41b8a8e9};
test_output[548] = '{32'h42409327};
/*############ DEBUG ############
test_input[4384:4391] = '{23.0824763469, 10.3340069663, -19.522597519, 34.4643682159, 21.897544802, -38.5446044098, 71.2261795345, -87.878169872};
test_label[548] = '{23.0824763469};
test_output[548] = '{48.1437031876};
############ END DEBUG ############*/
test_input[4392:4399] = '{32'hc2311e12, 32'h41a5f4c1, 32'h41840b65, 32'h42c36c9e, 32'hc283a1f0, 32'h4254ead9, 32'hc1453189, 32'hc2100e55};
test_label[549] = '{32'hc2311e12};
test_output[549] = '{32'h430dfdd3};
/*############ DEBUG ############
test_input[4392:4399] = '{-44.2793667339, 20.7445081313, 16.5055634108, 97.7121411397, -65.8162842692, 53.2293452271, -12.3245937914, -36.013996933};
test_label[549] = '{-44.2793667339};
test_output[549] = '{141.991507874};
############ END DEBUG ############*/
test_input[4400:4407] = '{32'h42942267, 32'h403e6dde, 32'hc2964d91, 32'hc28de99e, 32'h42117886, 32'h42b2c7fb, 32'h408f24f0, 32'h42916d21};
test_label[550] = '{32'hc2964d91};
test_output[550] = '{32'h43248ac6};
/*############ DEBUG ############
test_input[4400:4407] = '{74.0671946876, 2.97545580222, -75.151498963, -70.9562866747, 36.3676997917, 89.3905859381, 4.47325907454, 72.7131390703};
test_label[550] = '{-75.151498963};
test_output[550] = '{164.54208518};
############ END DEBUG ############*/
test_input[4408:4415] = '{32'hc2ac8c92, 32'hc29c10b9, 32'hc29d2eff, 32'hc09c736a, 32'h41785e16, 32'hc18862ab, 32'hc02bf741, 32'h41cc14f6};
test_label[551] = '{32'hc29d2eff};
test_output[551] = '{32'h42d03442};
/*############ DEBUG ############
test_input[4408:4415] = '{-86.2745490672, -78.0326607201, -78.5917882605, -4.88908877559, 15.5229705234, -17.0481786131, -2.68696612729, 25.5102343829};
test_label[551] = '{-78.5917882605};
test_output[551] = '{104.102068624};
############ END DEBUG ############*/
test_input[4416:4423] = '{32'h42c6c8c6, 32'hc2969d7f, 32'hc2827e20, 32'hbf81d78f, 32'h423d1544, 32'hc18fd3d7, 32'hc24a1f57, 32'h422341b6};
test_label[552] = '{32'hc2969d7f};
test_output[552] = '{32'h432eb323};
/*############ DEBUG ############
test_input[4416:4423] = '{99.3921367424, -75.3076122314, -65.2463406459, -1.01439081254, 47.2707673078, -17.9784366332, -50.5306057723, 40.8141719471};
test_label[552] = '{-75.3076122314};
test_output[552] = '{174.699748974};
############ END DEBUG ############*/
test_input[4424:4431] = '{32'hc2ab03ae, 32'hc1adb473, 32'hc267fadc, 32'h42136e35, 32'h42935903, 32'h42602d1a, 32'hc1e87d48, 32'hc0ff2c2a};
test_label[553] = '{32'h42935903};
test_output[553] = '{32'h32bd6f9d};
/*############ DEBUG ############
test_input[4424:4431] = '{-85.5071884178, -21.7131092315, -57.9949816801, 36.8576253991, 73.6738520012, 56.0440462468, -29.0611717094, -7.97414098648};
test_label[553] = '{73.6738520012};
test_output[553] = '{2.20532520235e-08};
############ END DEBUG ############*/
test_input[4432:4439] = '{32'hc2008923, 32'hc28f93ae, 32'hc2b00ada, 32'h4286398a, 32'h40ae1d8d, 32'h42841f7f, 32'hc2bf2046, 32'hc14bec40};
test_label[554] = '{32'hc2bf2046};
test_output[554] = '{32'h4322f9aa};
/*############ DEBUG ############
test_input[4432:4439] = '{-32.1339230193, -71.7884348939, -88.0211957908, 67.1123837406, 5.44110748783, 66.0615177432, -95.5630365376, -12.7451784428};
test_label[554] = '{-95.5630365376};
test_output[554] = '{162.975254342};
############ END DEBUG ############*/
test_input[4440:4447] = '{32'h4299afd7, 32'hc2496207, 32'h4259fae7, 32'hc1f3351a, 32'hc28dc0de, 32'hc27343ea, 32'hc10adac3, 32'hc27b06b8};
test_label[555] = '{32'h4259fae7};
test_output[555] = '{32'h41b2c990};
/*############ DEBUG ############
test_input[4440:4447] = '{76.8434385781, -50.345730458, 54.4950200631, -30.4009285477, -70.8766921731, -60.8163229469, -8.67840908933, -62.7565626413};
test_label[555] = '{54.4950200631};
test_output[555] = '{22.3484185152};
############ END DEBUG ############*/
test_input[4448:4455] = '{32'hc2b1bae8, 32'h41a56464, 32'h427f9a7d, 32'hc282a7ee, 32'hc1d363a1, 32'hc24884f7, 32'h4287cd98, 32'h41c90ac1};
test_label[556] = '{32'hc24884f7};
test_output[556] = '{32'h42ec195c};
/*############ DEBUG ############
test_input[4448:4455] = '{-88.8650542209, 20.6740189574, 63.9008688796, -65.3279865945, -26.4236470211, -50.1298469862, 67.9015476066, 25.1302507183};
test_label[556] = '{-50.1298469862};
test_output[556] = '{118.049532317};
############ END DEBUG ############*/
test_input[4456:4463] = '{32'hc268056a, 32'h4221bb14, 32'hc2b3c074, 32'h41556858, 32'hc2021a4a, 32'h4200e687, 32'h413d30ea, 32'h425ed2c1};
test_label[557] = '{32'h41556858};
test_output[557] = '{32'h422978ab};
/*############ DEBUG ############
test_input[4456:4463] = '{-58.0052884552, 40.4326920346, -89.8758816191, 13.3379749154, -32.5256714715, 32.2251260889, 11.8244418731, 55.705815905};
test_label[557] = '{13.3379749154};
test_output[557] = '{42.3678412224};
############ END DEBUG ############*/
test_input[4464:4471] = '{32'h4296808d, 32'h40817d31, 32'hc2a576fe, 32'h424bbeae, 32'hc2a2e032, 32'hc13f8659, 32'h42ae7ab2, 32'hc003fc2f};
test_label[558] = '{32'hc13f8659};
test_output[558] = '{32'h42c66b7e};
/*############ DEBUG ############
test_input[4464:4471] = '{75.2510763126, 4.04653198539, -82.7324082455, 50.9362107565, -81.4378813541, -11.9702996856, 87.2396360793, -2.06226710812};
test_label[558] = '{-11.9702996856};
test_output[558] = '{99.2099419798};
############ END DEBUG ############*/
test_input[4472:4479] = '{32'hc02bc8bb, 32'h42a8e56e, 32'h4233f7ee, 32'hc1613f96, 32'h4133c211, 32'h42650979, 32'h42c02d58, 32'hc22fb9ab};
test_label[559] = '{32'h4233f7ee};
test_output[559] = '{32'h424c62c4};
/*############ DEBUG ############
test_input[4472:4479] = '{-2.68412653724, 84.448103929, 44.9921179451, -14.0780242477, 11.2348793386, 57.2592522943, 96.0885590546, -43.9313171038};
test_label[559] = '{44.9921179451};
test_output[559] = '{51.0964499121};
############ END DEBUG ############*/
test_input[4480:4487] = '{32'h42938e9c, 32'hc21cdc81, 32'hc296bb05, 32'hc005cd70, 32'h42c2151f, 32'hc0adb259, 32'h42a82572, 32'h41305d11};
test_label[560] = '{32'h42c2151f};
test_output[560] = '{32'h361c9b8c};
/*############ DEBUG ############
test_input[4480:4487] = '{73.7785368455, -39.215337508, -75.3652760103, -2.09066385803, 97.0412522374, -5.42802108876, 84.0731362014, 11.022720849};
test_label[560] = '{97.0412522374};
test_output[560] = '{2.33363507484e-06};
############ END DEBUG ############*/
test_input[4488:4495] = '{32'hc2b40349, 32'hc2305a62, 32'hc22b3496, 32'hc1ec7b3b, 32'hc1d09295, 32'hc2c6278e, 32'h42260f04, 32'h421d137a};
test_label[561] = '{32'hc22b3496};
test_output[561] = '{32'h42a8d552};
/*############ DEBUG ############
test_input[4488:4495] = '{-90.0064159686, -44.0882633169, -42.8013518, -29.5601704246, -26.0715724791, -99.0772535909, 41.5146642305, 39.2690195871};
test_label[561] = '{-42.8013518};
test_output[561] = '{84.4166386894};
############ END DEBUG ############*/
test_input[4496:4503] = '{32'h427ca9fd, 32'hc18b4efd, 32'hc280fef5, 32'hc236c26e, 32'hc24d403c, 32'h42ac9b1f, 32'hc2855915, 32'h42a6a5db};
test_label[562] = '{32'hc18b4efd};
test_output[562] = '{32'h42cf8843};
/*############ DEBUG ############
test_input[4496:4503] = '{63.1660029126, -17.4135692499, -64.4979627101, -45.6898736587, -51.3127276012, 86.3029717123, -66.6739916225, 83.3239356994};
test_label[562] = '{-17.4135692499};
test_output[562] = '{103.76613254};
############ END DEBUG ############*/
test_input[4504:4511] = '{32'hc1368d86, 32'hc282ee66, 32'hc18e7826, 32'hc23c093a, 32'h42a0145c, 32'h426dd422, 32'hc0b40727, 32'hc24a9aec};
test_label[563] = '{32'hc282ee66};
test_output[563] = '{32'h43118161};
/*############ DEBUG ############
test_input[4504:4511] = '{-11.4095518503, -65.465622281, -17.8086659829, -47.0090116124, 80.0397654155, 59.4571605721, -5.62587330519, -50.6512899986};
test_label[563] = '{-65.465622281};
test_output[563] = '{145.505387698};
############ END DEBUG ############*/
test_input[4512:4519] = '{32'hc206314b, 32'h42c049b5, 32'hc28bfd1e, 32'hc2bc2eeb, 32'h42438b97, 32'hc25a8ac9, 32'h426bb8db, 32'hc1faa246};
test_label[564] = '{32'h426bb8db};
test_output[564] = '{32'h4214da90};
/*############ DEBUG ############
test_input[4512:4519] = '{-33.5481373061, 96.143962392, -69.9943660046, -94.091638518, 48.8863192307, -54.6355324955, 58.9305214757, -31.3292349065};
test_label[564] = '{58.9305214757};
test_output[564] = '{37.2134409163};
############ END DEBUG ############*/
test_input[4520:4527] = '{32'hc22847c3, 32'h4160d22a, 32'hc2178185, 32'h4122b024, 32'h3ff33da8, 32'hc268bbf7, 32'hc266f25d, 32'h41e40ced};
test_label[565] = '{32'h41e40ced};
test_output[565] = '{32'h3510880d};
/*############ DEBUG ############
test_input[4520:4527] = '{-42.0700799695, 14.0513093967, -37.8764857273, 10.1680031027, 1.90031905418, -58.183559263, -57.7366824234, 28.5063119354};
test_label[565] = '{28.5063119354};
test_output[565] = '{5.38421604699e-07};
############ END DEBUG ############*/
test_input[4528:4535] = '{32'h420d08fe, 32'hc1b21a97, 32'h429565a7, 32'h41ad38ea, 32'hc2292715, 32'hc0ebd777, 32'hc2945c33, 32'hc2978f46};
test_label[566] = '{32'h420d08fe};
test_output[566] = '{32'h421dc24f};
/*############ DEBUG ############
test_input[4528:4535] = '{35.2587826807, -22.2629831265, 74.6985374875, 21.6527901602, -42.288165129, -7.37005163198, -74.1800795703, -75.7798327585};
test_label[566] = '{35.2587826807};
test_output[566] = '{39.4397548068};
############ END DEBUG ############*/
test_input[4536:4543] = '{32'hc21e1117, 32'h414da8c9, 32'hc2bc8f35, 32'h40db2399, 32'h4286d7a9, 32'h427b99f0, 32'hc19666cc, 32'hc2b10e65};
test_label[567] = '{32'hc19666cc};
test_output[567] = '{32'h42ac76e6};
/*############ DEBUG ############
test_input[4536:4543] = '{-39.5166884618, 12.8537070746, -94.2796996148, 6.84809526677, 67.4212088582, 62.9003307141, -18.8001938798, -88.5281162083};
test_label[567] = '{-18.8001938798};
test_output[567] = '{86.2322234481};
############ END DEBUG ############*/
test_input[4544:4551] = '{32'h428da244, 32'hc266b4b3, 32'h4222b340, 32'h3f46d256, 32'h42ba747e, 32'hc1f0df24, 32'h4187b282, 32'hc27ca062};
test_label[568] = '{32'h428da244};
test_output[568] = '{32'h41b348e7};
/*############ DEBUG ############
test_input[4544:4551] = '{70.8169252687, -57.6764641386, 40.67504717, 0.776646981287, 93.2275212408, -30.1089547481, 16.962161906, -63.1566231558};
test_label[568] = '{70.8169252687};
test_output[568] = '{22.4105959723};
############ END DEBUG ############*/
test_input[4552:4559] = '{32'h426ccb5d, 32'hc21dbf99, 32'h42ac1bf6, 32'hc24e56d1, 32'hc2aa9fd6, 32'h429409e4, 32'hc23e61ee, 32'h42047928};
test_label[569] = '{32'hc24e56d1};
test_output[569] = '{32'h4309a3b0};
/*############ DEBUG ############
test_input[4552:4559] = '{59.1985980087, -39.4371071855, 86.0546115577, -51.5847826491, -85.312175972, 74.0193210036, -47.5956350285, 33.1183160608};
test_label[569] = '{-51.5847826491};
test_output[569] = '{137.639400138};
############ END DEBUG ############*/
test_input[4560:4567] = '{32'h41a0cf49, 32'hc2269ba1, 32'hc293f762, 32'h429b5b5b, 32'hc0868c2a, 32'hc1d24e8b, 32'h424adf46, 32'h41695d83};
test_label[570] = '{32'hc1d24e8b};
test_output[570] = '{32'h42cfeefe};
/*############ DEBUG ############
test_input[4560:4567] = '{20.1012129121, -41.6519813766, -73.9831697464, 77.6784288829, -4.20460983838, -26.2883501065, 50.7180413212, 14.5853298711};
test_label[570] = '{-26.2883501065};
test_output[570] = '{103.966778989};
############ END DEBUG ############*/
test_input[4568:4575] = '{32'hbf13ba27, 32'hc2a87639, 32'h41a7e9f0, 32'h42991dd6, 32'h41bacab7, 32'h42999a14, 32'h41dbf59d, 32'hc2c56550};
test_label[571] = '{32'hbf13ba27};
test_output[571] = '{32'h429bea10};
/*############ DEBUG ############
test_input[4568:4575] = '{-0.577059185278, -84.2309038581, 20.9892276974, 76.5582754092, 23.3489818142, 76.8009349002, 27.4949277752, -98.6978793717};
test_label[571] = '{-0.577059185278};
test_output[571] = '{77.957153986};
############ END DEBUG ############*/
test_input[4576:4583] = '{32'h42c01a0b, 32'h3e46945f, 32'hc2825baf, 32'hc2829e35, 32'h4255080b, 32'hc2c0b6a3, 32'h4294b29d, 32'h420def79};
test_label[572] = '{32'hc2829e35};
test_output[572] = '{32'h43215c20};
/*############ DEBUG ############
test_input[4576:4583] = '{96.0508614792, 0.193925371111, -65.1790682221, -65.3090008498, 53.2578538205, -96.3567121825, 74.3488563762, 35.4838612347};
test_label[572] = '{-65.3090008498};
test_output[572] = '{161.359862329};
############ END DEBUG ############*/
test_input[4584:4591] = '{32'hc2544118, 32'h419a98a6, 32'h425f6b39, 32'h429ee282, 32'h426fe917, 32'hc1c71a86, 32'hc28b3467, 32'h42a957b9};
test_label[573] = '{32'hc28b3467};
test_output[573] = '{32'h431a476f};
/*############ DEBUG ############
test_input[4584:4591] = '{-53.0635665396, 19.3245345511, 55.8547077249, 79.4423953415, 59.977628254, -24.8879502224, -69.6023520341, 84.6713365428};
test_label[573] = '{-69.6023520341};
test_output[573] = '{154.279033464};
############ END DEBUG ############*/
test_input[4592:4599] = '{32'h425e0149, 32'hc275d1e2, 32'hc29df08f, 32'h4217f1e1, 32'hc2c7733f, 32'h4234405b, 32'hc2991a66, 32'h4238614f};
test_label[574] = '{32'hc2c7733f};
test_output[574] = '{32'h431b39f9};
/*############ DEBUG ############
test_input[4592:4599] = '{55.5012551471, -61.4549633289, -78.9698431108, 37.986211467, -99.7250911953, 45.0628466546, -76.5515595128, 46.095026913};
test_label[574] = '{-99.7250911953};
test_output[574] = '{155.226457857};
############ END DEBUG ############*/
test_input[4600:4607] = '{32'hc209f643, 32'hc17b72b9, 32'h40c0578a, 32'hc2c49d26, 32'hc2a477d7, 32'h42282e66, 32'h41d3f117, 32'h42c7459b};
test_label[575] = '{32'h42282e66};
test_output[575] = '{32'h42665cd0};
/*############ DEBUG ############
test_input[4600:4607] = '{-34.4904902701, -15.7155081533, 6.01068596794, -98.3069281804, -82.2340626909, 42.04531072, 26.4927203053, 99.6359491037};
test_label[575] = '{42.04531072};
test_output[575] = '{57.5906383837};
############ END DEBUG ############*/
test_input[4608:4615] = '{32'h42c01791, 32'hc22109da, 32'hc19d19f6, 32'hc1e0a3df, 32'h41e3df82, 32'hc24833f0, 32'h428dd286, 32'hc0cb181d};
test_label[576] = '{32'hc24833f0};
test_output[576] = '{32'h431218c5};
/*############ DEBUG ############
test_input[4608:4615] = '{96.0460308335, -40.2596213773, -19.6376753796, -28.0800146607, 28.4841340919, -50.0507184912, 70.9111800722, -6.34669365149};
test_label[576] = '{-50.0507184912};
test_output[576] = '{146.096749325};
############ END DEBUG ############*/
test_input[4616:4623] = '{32'hc2863b7e, 32'hc2993e6e, 32'hc2823e82, 32'hc21d7b13, 32'hc2c414c6, 32'hc17369b2, 32'hc28ca2ae, 32'hc108d531};
test_label[577] = '{32'hc28ca2ae};
test_output[577] = '{32'h4277115f};
/*############ DEBUG ############
test_input[4616:4623] = '{-67.1161944113, -76.6219332324, -65.1220886876, -39.370190127, -98.0405694766, -15.2133040505, -70.3177336872, -8.55204888977};
test_label[577] = '{-70.3177336872};
test_output[577] = '{61.7669635188};
############ END DEBUG ############*/
test_input[4624:4631] = '{32'hc26ec875, 32'h412c6ae2, 32'hc1a2befe, 32'h4231c2d2, 32'h42433a07, 32'hc01082c7, 32'hc203317e, 32'h41ebfebb};
test_label[578] = '{32'h412c6ae2};
test_output[578] = '{32'h42182c3a};
/*############ DEBUG ############
test_input[4624:4631] = '{-59.6957575645, 10.7760943545, -20.343257541, 44.4402556853, 48.8066688025, -2.25798198093, -32.7983324379, 29.4993806541};
test_label[578] = '{10.7760943545};
test_output[578] = '{38.0431912254};
############ END DEBUG ############*/
test_input[4632:4639] = '{32'hc1a9c320, 32'hc1dbd260, 32'hc29c4090, 32'hc1c6fe3b, 32'hc2a29382, 32'h406a9045, 32'h42c2b296, 32'h42b184a3};
test_label[579] = '{32'hc29c4090};
test_output[579] = '{32'h432f799f};
/*############ DEBUG ############
test_input[4632:4639] = '{-21.220275157, -27.4777215306, -78.1260951519, -24.8741355263, -81.2881005242, 3.66505542864, 97.3487978213, 88.7590540288};
test_label[579] = '{-78.1260951519};
test_output[579] = '{175.47507896};
############ END DEBUG ############*/
test_input[4640:4647] = '{32'h423534a7, 32'hc2b3e2b9, 32'h42ba8f4d, 32'h419f873e, 32'hc1ad0c30, 32'h4294d970, 32'h410e6681, 32'h41b0e7f7};
test_label[580] = '{32'h42ba8f4d};
test_output[580] = '{32'h31de8102};
/*############ DEBUG ############
test_input[4640:4647] = '{45.3014201115, -89.9428200484, 93.2798859366, 19.941036199, -21.6309502772, 74.4246794158, 8.90002579817, 22.1132634755};
test_label[580] = '{93.2798859366};
test_output[580] = '{6.47571676158e-09};
############ END DEBUG ############*/
test_input[4648:4655] = '{32'h428da8ca, 32'h42982b86, 32'hc089ed6a, 32'h42af19f1, 32'h42990387, 32'h42938573, 32'hc2af83ba, 32'h42acedbe};
test_label[581] = '{32'hc2af83ba};
test_output[581] = '{32'h432f9947};
/*############ DEBUG ############
test_input[4648:4655] = '{70.8296632124, 76.0850081814, -4.31023125688, 87.5506679233, 76.5068882692, 73.7606401617, -87.7572776442, 86.4643380616};
test_label[581] = '{-87.7572776442};
test_output[581] = '{175.598733018};
############ END DEBUG ############*/
test_input[4656:4663] = '{32'h42b13bfc, 32'hc1df813f, 32'h4034226a, 32'h42a24094, 32'hc29c57e1, 32'hc252ba8c, 32'h4287f9dc, 32'h42909983};
test_label[582] = '{32'h42909983};
test_output[582] = '{32'h41828b0c};
/*############ DEBUG ############
test_input[4656:4663] = '{88.6171592553, -27.9381092495, 2.81460040248, 81.1261258968, -78.1716394874, -52.6821738294, 67.9880067006, 72.299824059};
test_label[582] = '{72.299824059};
test_output[582] = '{16.3178931897};
############ END DEBUG ############*/
test_input[4664:4671] = '{32'h42c44291, 32'hc2ae1ee6, 32'h42b8710f, 32'h4229f39f, 32'hc22ead0e, 32'hc18ee071, 32'h420bd43b, 32'hc2bcfc1e};
test_label[583] = '{32'hc2bcfc1e};
test_output[583] = '{32'h4340a009};
/*############ DEBUG ############
test_input[4664:4671] = '{98.1300121977, -87.0603474618, 92.2208139989, 42.4879111356, -43.6689994883, -17.859591182, 34.9572580363, -94.4924192719};
test_label[583] = '{-94.4924192719};
test_output[583] = '{192.625142155};
############ END DEBUG ############*/
test_input[4672:4679] = '{32'h4278bb74, 32'hc1b71003, 32'hc07fd6ee, 32'h421ced78, 32'hc1c460a2, 32'hc25f7b59, 32'h425eb6c0, 32'hc18544dd};
test_label[584] = '{32'hc1b71003};
test_output[584] = '{32'h42aa227f};
/*############ DEBUG ############
test_input[4672:4679] = '{62.183060756, -22.8828182618, -3.99749334602, 39.2319012439, -24.5471833893, -55.8704572332, 55.6784653533, -16.6586252782};
test_label[584] = '{-22.8828182618};
test_output[584] = '{85.0673744453};
############ END DEBUG ############*/
test_input[4680:4687] = '{32'hc219cafb, 32'hc27b3658, 32'h40a8e9eb, 32'hc250b254, 32'hc28b2161, 32'hc2831564, 32'h4198de5e, 32'h40f33bcf};
test_label[585] = '{32'hc2831564};
test_output[585] = '{32'h42a94cfd};
/*############ DEBUG ############
test_input[4680:4687] = '{-38.448223095, -62.8030692823, 5.27855428726, -52.1741485826, -69.5651943106, -65.5417809135, 19.1085771224, 7.60105102204};
test_label[585] = '{-65.5417809135};
test_output[585] = '{84.6503690756};
############ END DEBUG ############*/
test_input[4688:4695] = '{32'h42809ba4, 32'hc1dda16c, 32'hc1273452, 32'h41b76a5d, 32'h427a53e9, 32'h40e387c1, 32'h424157aa, 32'hc2aab07a};
test_label[586] = '{32'h40e387c1};
test_output[586] = '{32'h42656eac};
/*############ DEBUG ############
test_input[4688:4695] = '{64.3039869426, -27.7038189876, -10.4502732577, 22.926934633, 62.5819426831, 7.11032137225, 48.3356106878, -85.344678739};
test_label[586] = '{7.11032137225};
test_output[586] = '{57.3580781989};
############ END DEBUG ############*/
test_input[4696:4703] = '{32'h42c38ec9, 32'hc26aae9f, 32'h428b0279, 32'h42b39f15, 32'h4144c3ce, 32'h42035274, 32'hc29c60a4, 32'hc0e555b8};
test_label[587] = '{32'h4144c3ce};
test_output[587] = '{32'h42aaf67d};
/*############ DEBUG ############
test_input[4696:4703] = '{97.7788806065, -58.6705293597, 69.5048318194, 89.8107078643, 12.2978038063, 32.8305219401, -78.1887490591, -7.16671356651};
test_label[587] = '{12.2978038063};
test_output[587] = '{85.4814230515};
############ END DEBUG ############*/
test_input[4704:4711] = '{32'h429abb72, 32'hc1f62a65, 32'h4297772d, 32'hc282538d, 32'hc22ae9ed, 32'hc152398a, 32'h426a7702, 32'hc1fe854c};
test_label[588] = '{32'hc22ae9ed};
test_output[588] = '{32'h42f08bbd};
/*############ DEBUG ############
test_input[4704:4711] = '{77.366107639, -30.7707004516, 75.7327667234, -65.163188187, -42.7284441619, -13.139047317, 58.6162171458, -31.815086416};
test_label[588] = '{-42.7284441619};
test_output[588] = '{120.272928997};
############ END DEBUG ############*/
test_input[4712:4719] = '{32'h42bd100f, 32'hc2b4af84, 32'hc22a6e42, 32'hc222303a, 32'hc2bbe41e, 32'h41aa6009, 32'hc1fc200b, 32'h42662d65};
test_label[589] = '{32'hc2bbe41e};
test_output[589] = '{32'h433c7a16};
/*############ DEBUG ############
test_input[4712:4719] = '{94.5313649557, -90.3428076106, -42.6076718728, -40.5470957312, -93.9455397217, 21.2968924865, -31.515645625, 57.5443322408};
test_label[589] = '{-93.9455397217};
test_output[589] = '{188.476904677};
############ END DEBUG ############*/
test_input[4720:4727] = '{32'hc226c679, 32'hc1fc9344, 32'h422faef7, 32'h422b59f7, 32'h42ba5204, 32'h4234f093, 32'h42bb31a3, 32'h429ab75c};
test_label[590] = '{32'h42bb31a3};
test_output[590] = '{32'h3eff31b6};
/*############ DEBUG ############
test_input[4720:4727] = '{-41.6938217871, -31.5719079361, 43.9208635449, 42.8378551497, 93.1601904238, 45.2349362007, 93.5969475123, 77.3581209133};
test_label[590] = '{93.5969475123};
test_output[590] = '{0.498426138679};
############ END DEBUG ############*/
test_input[4728:4735] = '{32'h41a8c3b4, 32'hc2021eed, 32'hc1cf0f8f, 32'h42832b7e, 32'hc20673a7, 32'hc27bba35, 32'hc0c652d7, 32'hc07cd7b1};
test_label[591] = '{32'hc20673a7};
test_output[591] = '{32'h42c66552};
/*############ DEBUG ############
test_input[4728:4735] = '{21.0955575952, -32.5302020596, -25.8825960399, 65.5849456489, -33.6129423028, -62.9318426142, -6.19761224622, -3.95066479461};
test_label[591] = '{-33.6129423028};
test_output[591] = '{99.1978879517};
############ END DEBUG ############*/
test_input[4736:4743] = '{32'h42b25e6d, 32'h420a51c3, 32'hc28d7953, 32'h42b6c7fa, 32'hc212f62b, 32'hc288970e, 32'h42c6b138, 32'h426b3235};
test_label[592] = '{32'h420a51c3};
test_output[592] = '{32'h4281888a};
/*############ DEBUG ############
test_input[4736:4743] = '{89.1844239554, 34.5798470656, -70.7369644388, 91.3905791409, -36.7403966094, -68.2950310508, 99.346133138, 58.7990294831};
test_label[592] = '{34.5798470656};
test_output[592] = '{64.7666753268};
############ END DEBUG ############*/
test_input[4744:4751] = '{32'h4270c199, 32'hc20f158e, 32'hc230108c, 32'h42bb0dd5, 32'hc2987f70, 32'h3f95c8a0, 32'hc26cc732, 32'hc2ae44ce};
test_label[593] = '{32'h3f95c8a0};
test_output[593] = '{32'h42b8b6b2};
/*############ DEBUG ############
test_input[4744:4751] = '{60.1890609999, -35.771050588, -44.016159748, 93.5270134341, -76.2488986259, 1.17018512606, -59.1945277759, -87.1343847109};
test_label[593] = '{1.17018512606};
test_output[593] = '{92.3568283081};
############ END DEBUG ############*/
test_input[4752:4759] = '{32'hc2a10f64, 32'hc25006e6, 32'h4264ac9b, 32'h4292030c, 32'h42c7e58b, 32'hc20f3fe4, 32'hc2432874, 32'hc2bd4651};
test_label[594] = '{32'hc25006e6};
test_output[594] = '{32'h4317f47f};
/*############ DEBUG ############
test_input[4752:4759] = '{-80.530060417, -52.0067354912, 57.1685586409, 73.0059515414, 99.9483238776, -35.8123950844, -48.7895054561, -94.6373384085};
test_label[594] = '{-52.0067354912};
test_output[594] = '{151.955059369};
############ END DEBUG ############*/
test_input[4760:4767] = '{32'hc28a51ca, 32'h421959cd, 32'hc01b48e5, 32'hc29e98ca, 32'h428ab5f7, 32'h424aad8d, 32'h42c57f51, 32'hc275bad3};
test_label[595] = '{32'h424aad8d};
test_output[595] = '{32'h42405116};
/*############ DEBUG ############
test_input[4760:4767] = '{-69.1597445283, 38.3376958911, -2.42632408946, -79.2984189065, 69.3554029327, 50.6694819629, 98.7486672255, -61.43244667};
test_label[595] = '{50.6694819629};
test_output[595] = '{48.0791852626};
############ END DEBUG ############*/
test_input[4768:4775] = '{32'hc2c4965a, 32'h4236f814, 32'hc29a3498, 32'hc2685fc8, 32'hc19cb83e, 32'hc182f270, 32'hc282104d, 32'h425e2b92};
test_label[596] = '{32'hc29a3498};
test_output[596] = '{32'h4304a534};
/*############ DEBUG ############
test_input[4768:4775] = '{-98.293651922, 45.7422649923, -77.1027259215, -58.0935380469, -19.5899628698, -16.3683775108, -65.03183374, 55.5425492224};
test_label[596] = '{-77.1027259215};
test_output[596] = '{132.645330578};
############ END DEBUG ############*/
test_input[4776:4783] = '{32'hc2894096, 32'hc26a6989, 32'h42aa39f0, 32'hc17f8461, 32'hc1bde6d7, 32'h42817be0, 32'hc0dc83c1, 32'h42a23100};
test_label[597] = '{32'h42a23100};
test_output[597] = '{32'h4081211b};
/*############ DEBUG ############
test_input[4776:4783] = '{-68.62614334, -58.6030608525, 85.1131579237, -15.9698189519, -23.7377141664, 64.7419466794, -6.89108312706, 81.0957053438};
test_label[597] = '{81.0957053438};
test_output[597] = '{4.03529127835};
############ END DEBUG ############*/
test_input[4784:4791] = '{32'hc0c51249, 32'h41baee43, 32'h4260bb0c, 32'h42449db3, 32'hc2b74d87, 32'h4203a47c, 32'hc17ac050, 32'hc297a0c0};
test_label[598] = '{32'hc297a0c0};
test_output[598] = '{32'h4303ff5d};
/*############ DEBUG ############
test_input[4784:4791] = '{-6.1584818823, 23.3663389323, 56.1826638349, 49.1540024396, -91.6514193234, 32.9106284363, -15.6719510215, -75.8139625831};
test_label[598] = '{-75.8139625831};
test_output[598] = '{131.997512143};
############ END DEBUG ############*/
test_input[4792:4799] = '{32'h40f4c561, 32'h42a9cbde, 32'h4220cdfd, 32'hc0af7d4a, 32'hc2508251, 32'h40247c69, 32'h4125c31d, 32'hc2b49d3e};
test_label[599] = '{32'hc2508251};
test_output[599] = '{32'h43090683};
/*############ DEBUG ############
test_input[4792:4799] = '{7.6490939322, 84.8981787396, 40.2011599256, -5.48404401662, -52.1272634775, 2.5700934833, 10.3601350327, -90.307109876};
test_label[599] = '{-52.1272634775};
test_output[599] = '{137.025442217};
############ END DEBUG ############*/
test_input[4800:4807] = '{32'h4239359c, 32'hc028897c, 32'h42b3c095, 32'h41e779ab, 32'h41836809, 32'h429b9e48, 32'hc234507e, 32'hc2a0c498};
test_label[600] = '{32'h4239359c};
test_output[600] = '{32'h422e4b90};
/*############ DEBUG ############
test_input[4800:4807] = '{46.3023532801, -2.63339132163, 89.8761374782, 28.9344082943, 16.425799172, 77.8091414356, -45.0786054374, -80.3839712817};
test_label[600] = '{46.3023532801};
test_output[600] = '{43.5737899442};
############ END DEBUG ############*/
test_input[4808:4815] = '{32'hbe19cc20, 32'hc2a89d47, 32'hc27e8095, 32'hc19f2316, 32'h421ddd1e, 32'hc180e78f, 32'hbfc5a0a0, 32'h41fc10b8};
test_label[601] = '{32'hc2a89d47};
test_output[601] = '{32'h42f78c04};
/*############ DEBUG ############
test_input[4808:4815] = '{-0.150192740636, -84.3071844703, -63.6255680568, -19.8921311278, 39.4659348368, -16.1130652104, -1.54396438953, 31.5081632264};
test_label[601] = '{-84.3071844703};
test_output[601] = '{123.773469178};
############ END DEBUG ############*/
test_input[4816:4823] = '{32'hc27f071f, 32'h4254eca2, 32'h42889c73, 32'h404b2b05, 32'h41cb0fe1, 32'h4259ff4a, 32'h420bdcf4, 32'hc29e518e};
test_label[602] = '{32'hc27f071f};
test_output[602] = '{32'h43041001};
/*############ DEBUG ############
test_input[4816:4823] = '{-63.7569539217, 53.2310864812, 68.3055640588, 3.17450073526, 25.3827534202, 54.4993073132, 34.9657730796, -79.1592847661};
test_label[602] = '{-63.7569539217};
test_output[602] = '{132.062519274};
############ END DEBUG ############*/
test_input[4824:4831] = '{32'h4036e6c2, 32'hc2267211, 32'h420cf7b3, 32'h41f4e526, 32'hc1a6cc27, 32'hc20c97ae, 32'hc0a652bf, 32'hc28a7bec};
test_label[603] = '{32'h4036e6c2};
test_output[603] = '{32'h42019338};
/*############ DEBUG ############
test_input[4824:4831] = '{2.85783436429, -41.6113941936, 35.2418947878, 30.6118882204, -20.8496828259, -35.1481258832, -5.19760079959, -69.2420355646};
test_label[603] = '{2.85783436429};
test_output[603] = '{32.3937678486};
############ END DEBUG ############*/
test_input[4832:4839] = '{32'h427d0b48, 32'h428673c8, 32'h42c5519b, 32'h42110cb0, 32'h42b1564c, 32'h42b987ba, 32'h42b14bc4, 32'h41b51ade};
test_label[604] = '{32'h427d0b48};
test_output[604] = '{32'h420d9ad6};
/*############ DEBUG ############
test_input[4832:4839] = '{63.261017854, 67.2261377574, 98.6593843426, 36.2623896796, 88.6685489976, 92.765093553, 88.6479762968, 22.6381184111};
test_label[604] = '{63.261017854};
test_output[604] = '{35.4012082794};
############ END DEBUG ############*/
test_input[4840:4847] = '{32'hc179ff37, 32'h4219cc96, 32'h42ad3455, 32'h423c05ba, 32'hc29af46e, 32'hc19af52a, 32'h42ad1862, 32'h428c4448};
test_label[605] = '{32'hc19af52a};
test_output[605] = '{32'h42d546bb};
/*############ DEBUG ############
test_input[4840:4847] = '{-15.6248087431, 38.4497908437, 86.6022098271, 47.0055934079, -77.4774052188, -19.3697096767, 86.547623961, 70.1333636426};
test_label[605] = '{-19.3697096767};
test_output[605] = '{106.638146193};
############ END DEBUG ############*/
test_input[4848:4855] = '{32'hc11c4fd3, 32'hc2717175, 32'hc2afa0c2, 32'hc2bf239e, 32'hc11f0b5a, 32'hc162669a, 32'h41539569, 32'h42703883};
test_label[606] = '{32'h41539569};
test_output[606] = '{32'h423b5329};
/*############ DEBUG ############
test_input[4848:4855] = '{-9.76948816469, -60.3607983529, -87.813980732, -95.569561597, -9.94027138688, -14.1500494429, 13.2239770159, 60.0551879504};
test_label[606] = '{13.2239770159};
test_output[606] = '{46.8312109345};
############ END DEBUG ############*/
test_input[4856:4863] = '{32'hc2a3e92e, 32'hc24582d8, 32'hc26a5014, 32'h42c00ef2, 32'h4248cb72, 32'hbfa7423c, 32'hc291e51e, 32'h41d74aa7};
test_label[607] = '{32'hbfa7423c};
test_output[607] = '{32'h42c2abfb};
/*############ DEBUG ############
test_input[4856:4863] = '{-81.9554299798, -49.3777765875, -58.5782031088, 96.0291917975, 50.1986756076, -1.30670880505, -72.9474964426, 26.9114521706};
test_label[607] = '{-1.30670880505};
test_output[607] = '{97.3359006025};
############ END DEBUG ############*/
test_input[4864:4871] = '{32'hc20e3192, 32'hc1911901, 32'h42a1b31e, 32'h4167e3f0, 32'hc14042be, 32'h4274a4e6, 32'h41ef8635, 32'hc1c34961};
test_label[608] = '{32'hc1911901};
test_output[608] = '{32'h42c5f95e};
/*############ DEBUG ############
test_input[4864:4871] = '{-35.5484078358, -18.137208179, 80.8498393206, 14.4931484756, -12.0162947545, 61.1610340514, 29.9405312015, -24.4108302365};
test_label[608] = '{-18.137208179};
test_output[608] = '{98.9870475023};
############ END DEBUG ############*/
test_input[4872:4879] = '{32'h4298823e, 32'hc2a7e24e, 32'h42c3283d, 32'h42a530fb, 32'hc2b7385f, 32'hc2225993, 32'hc0f51af1, 32'hc1ac4c22};
test_label[609] = '{32'hc2b7385f};
test_output[609] = '{32'h433d304e};
/*############ DEBUG ############
test_input[4872:4879] = '{76.25438256, -83.9419980583, 97.5785936611, 82.5956645983, -91.6101013778, -40.5874741847, -7.65953854881, -21.5371744749};
test_label[609] = '{-91.6101013778};
test_output[609] = '{189.188695351};
############ END DEBUG ############*/
test_input[4880:4887] = '{32'h4143ae8e, 32'h41e715f8, 32'h4245a60c, 32'h41d5f023, 32'h42ae97a4, 32'hc2b85275, 32'hc28fc9a3, 32'hc2a1dd25};
test_label[610] = '{32'hc28fc9a3};
test_output[610] = '{32'h431f30a3};
/*############ DEBUG ############
test_input[4880:4887] = '{12.2301159926, 28.8857261804, 49.4121538828, 26.7422533352, 87.2961692816, -92.1610505756, -71.8938230678, -80.9319261812};
test_label[610] = '{-71.8938230678};
test_output[610] = '{159.189992349};
############ END DEBUG ############*/
test_input[4888:4895] = '{32'hc25c5710, 32'h42848d98, 32'h42c2fca7, 32'h3f95f82f, 32'h42ad9072, 32'h421b6595, 32'hc2a0bf28, 32'hc1e81573};
test_label[611] = '{32'hc25c5710};
test_output[611] = '{32'h43189419};
/*############ DEBUG ############
test_input[4888:4895] = '{-55.0850223332, 66.276547731, 97.4934615346, 1.17163646032, 86.7821220595, 38.8492012284, -80.3733483382, -29.0104738611};
test_label[611] = '{-55.0850223332};
test_output[611] = '{152.578506158};
############ END DEBUG ############*/
test_input[4896:4903] = '{32'hc24c3a25, 32'hc2138376, 32'hc26f6469, 32'h421c1462, 32'hc26a6070, 32'h41a13028, 32'hc27642ec, 32'hc2a8712c};
test_label[612] = '{32'h41a13028};
test_output[612] = '{32'h4196f89c};
/*############ DEBUG ############
test_input[4896:4903] = '{-51.0567833546, -36.8783780478, -59.8480564587, 39.0199065693, -58.5941783228, 20.1485145721, -61.5653525841, -84.2210422397};
test_label[612] = '{20.1485145721};
test_output[612] = '{18.8713920037};
############ END DEBUG ############*/
test_input[4904:4911] = '{32'h423ddf14, 32'h42c204f2, 32'h42af5176, 32'hc0ca1974, 32'h42aa59c4, 32'hc2164efc, 32'h41122a19, 32'h423c1341};
test_label[613] = '{32'hc0ca1974};
test_output[613] = '{32'h42cea696};
/*############ DEBUG ############
test_input[4904:4911] = '{47.4678505213, 97.0096601313, 87.6591052861, -6.31560701128, 85.175327082, -37.577132862, 9.13527802731, 47.0188040796};
test_label[613] = '{-6.31560701128};
test_output[613] = '{103.325361307};
############ END DEBUG ############*/
test_input[4912:4919] = '{32'h42530f3c, 32'h42173099, 32'h421a688d, 32'h4297b47f, 32'hc26f2b41, 32'h4168a867, 32'h40a6ce23, 32'hc1d6c92e};
test_label[614] = '{32'h4297b47f};
test_output[614] = '{32'h2eceb920};
/*############ DEBUG ############
test_input[4912:4919] = '{52.7648780443, 37.7974567909, 38.6021008888, 75.8525326306, -59.7922414978, 14.5411134881, 5.21266309363, -26.8482314391};
test_label[614] = '{75.8525326306};
test_output[614] = '{9.40068023469e-11};
############ END DEBUG ############*/
test_input[4920:4927] = '{32'hc17c0074, 32'hc29d3add, 32'h4187d54b, 32'h4263cb1d, 32'h41b0d384, 32'hc196b9de, 32'hc25de6fb, 32'hc2b45851};
test_label[615] = '{32'h41b0d384};
test_output[615] = '{32'h420b615b};
/*############ DEBUG ############
test_input[4920:4927] = '{-15.7501104021, -78.6149708392, 16.9791476462, 56.9483531197, 22.10327839, -18.8407545462, -55.4755657224, -90.1724963739};
test_label[615] = '{22.10327839};
test_output[615] = '{34.8450747297};
############ END DEBUG ############*/
test_input[4928:4935] = '{32'h421ad7a9, 32'hc0bb26e7, 32'h416ba537, 32'h42945257, 32'h42a807ed, 32'h4104b23e, 32'hc2c1ddcf, 32'hc2800d28};
test_label[616] = '{32'hc0bb26e7};
test_output[616] = '{32'h42b3ba63};
/*############ DEBUG ############
test_input[4928:4935] = '{38.7106045857, -5.84849890709, 14.7278354519, 74.1608213266, 84.0154821947, 8.29351661717, -96.9332180435, -64.0256944418};
test_label[616] = '{-5.84849890709};
test_output[616] = '{89.8640336023};
############ END DEBUG ############*/
test_input[4936:4943] = '{32'h40cd7470, 32'hc142c6e0, 32'hbfbf1827, 32'hc116a604, 32'h425195e3, 32'h4267ef60, 32'h4247bff6, 32'hc225d84c};
test_label[617] = '{32'h40cd7470};
test_output[617] = '{32'h424e44f9};
/*############ DEBUG ############
test_input[4936:4943] = '{6.42046349285, -12.1735538398, -1.4929246167, -9.41553106938, 52.3963755857, 57.9837642858, 49.937462412, -41.4612286205};
test_label[617] = '{6.42046349285};
test_output[617] = '{51.567357631};
############ END DEBUG ############*/
test_input[4944:4951] = '{32'hc2387371, 32'h42781a9d, 32'h429828cd, 32'h429272ba, 32'hc2561f2e, 32'hbf88ef06, 32'hc072a753, 32'h411de59c};
test_label[618] = '{32'hbf88ef06};
test_output[618] = '{32'h429a692b};
/*############ DEBUG ############
test_input[4944:4951] = '{-46.1127359722, 62.0259881535, 76.0796870687, 73.224079097, -53.5304504289, -1.06979440314, -3.7914626795, 9.86855667889};
test_label[618] = '{-1.06979440314};
test_output[618] = '{77.2054095551};
############ END DEBUG ############*/
test_input[4952:4959] = '{32'hc068e96e, 32'h42372739, 32'h42474b60, 32'hc2a3de65, 32'hc1ee9a8a, 32'h421357d0, 32'hc2312110, 32'h4233b0a0};
test_label[619] = '{32'hc068e96e};
test_output[619] = '{32'h4255f35f};
/*############ DEBUG ############
test_input[4952:4959] = '{-3.6392474606, 45.7883049971, 49.8236083591, -81.9343666404, -29.8254579139, 36.83575398, -44.2822866504, 44.9224840939};
test_label[619] = '{-3.6392474606};
test_output[619] = '{53.4876662981};
############ END DEBUG ############*/
test_input[4960:4967] = '{32'hc2b1607e, 32'h42c32114, 32'h41c399c9, 32'h428012bb, 32'hc29511ce, 32'h4283b694, 32'h420c9281, 32'hc1ab2dba};
test_label[620] = '{32'hc2b1607e};
test_output[620] = '{32'h433a40c9};
/*############ DEBUG ############
test_input[4960:4967] = '{-88.6884592069, 97.5646029991, 24.4500898321, 64.0365796847, -74.5347716454, 65.8565970632, 35.1430707575, -21.3973275845};
test_label[620] = '{-88.6884592069};
test_output[620] = '{186.253062206};
############ END DEBUG ############*/
test_input[4968:4975] = '{32'hc1c3d7d9, 32'h429a268c, 32'hc2c2ccdb, 32'hc29575a8, 32'h42c7df3c, 32'hc09b132a, 32'h41d65f60, 32'h422e26ce};
test_label[621] = '{32'hc1c3d7d9};
test_output[621] = '{32'h42f8d532};
/*############ DEBUG ############
test_input[4968:4975] = '{-24.4803940393, 77.0752856408, -97.4001059398, -74.7297970571, 99.9360022098, -4.8460894239, 26.7965704593, 43.5378936834};
test_label[621] = '{-24.4803940393};
test_output[621] = '{124.416396249};
############ END DEBUG ############*/
test_input[4976:4983] = '{32'hc2bfde51, 32'h42983750, 32'h41d18e36, 32'hc19bc19b, 32'h42ab1718, 32'hc21e0aae, 32'h412dbee1, 32'h4213d936};
test_label[622] = '{32'h42ab1718};
test_output[622] = '{32'h38a72a04};
/*############ DEBUG ############
test_input[4976:4983] = '{-95.9342122678, 76.1080317809, 26.1944385658, -19.4695344221, 85.5451066095, -39.5104299618, 10.8591015038, 36.9621191919};
test_label[622] = '{85.5451066095};
test_output[622] = '{7.97100658068e-05};
############ END DEBUG ############*/
test_input[4984:4991] = '{32'hc0546295, 32'hc24b35a6, 32'hc29e7f1b, 32'h425b08d5, 32'h42097fa5, 32'hc2843597, 32'h419afc67, 32'h4181b4c3};
test_label[623] = '{32'h4181b4c3};
test_output[623] = '{32'h421a2e73};
/*############ DEBUG ############
test_input[4984:4991] = '{-3.31851704188, -50.8023921179, -79.2482514837, 54.7586243808, 34.3746541665, -66.1046660107, 19.3732425343, 16.2132630265};
test_label[623] = '{16.2132630265};
test_output[623] = '{38.5453613557};
############ END DEBUG ############*/
test_input[4992:4999] = '{32'hc2ab0b62, 32'hc1c6d2dd, 32'h420cd4f9, 32'hc2660d07, 32'hc2c2b0a7, 32'hc02f2576, 32'h425b459e, 32'h42933c21};
test_label[624] = '{32'hc2c2b0a7};
test_output[624] = '{32'h432af664};
/*############ DEBUG ############
test_input[4992:4999] = '{-85.52223567, -24.8529609314, 35.2079824234, -57.5127214255, -97.3450261372, -2.73666139851, 54.8179854989, 73.6174381668};
test_label[624] = '{-97.3450261372};
test_output[624] = '{170.962464311};
############ END DEBUG ############*/
test_input[5000:5007] = '{32'h42b71b04, 32'h42433267, 32'h429eeeb9, 32'hc21c7aed, 32'h428ecb00, 32'hc1a792cb, 32'hc278923c, 32'h42a5c9e0};
test_label[625] = '{32'h42433267};
test_output[625] = '{32'h422b03d0};
/*############ DEBUG ############
test_input[5000:5007] = '{91.5527649937, 48.7992211611, 79.4662538365, -39.1200462353, 71.3964809967, -20.9466767987, -62.1428078294, 82.8942891837};
test_label[625] = '{48.7992211611};
test_output[625] = '{42.753723102};
############ END DEBUG ############*/
test_input[5008:5015] = '{32'h4290b95d, 32'h4040fa82, 32'h41c4e3d4, 32'hc21ced01, 32'hc295aeda, 32'h423039c0, 32'h40e60d60, 32'h42139c59};
test_label[626] = '{32'hc21ced01};
test_output[626] = '{32'h42df2fde};
/*############ DEBUG ############
test_input[5008:5015] = '{72.3620388354, 3.01528974338, 24.611243511, -39.2314484225, -74.8415050259, 44.0563973791, 7.18913261679, 36.9026820805};
test_label[626] = '{-39.2314484225};
test_output[626] = '{111.593487258};
############ END DEBUG ############*/
test_input[5016:5023] = '{32'h42349ccb, 32'h4283f260, 32'h427e4b69, 32'h4203c6e4, 32'hc2ad4674, 32'h42414731, 32'hc25843ce, 32'hc294c46f};
test_label[627] = '{32'hc25843ce};
test_output[627] = '{32'h42f040bf};
/*############ DEBUG ############
test_input[5016:5023] = '{45.1531189471, 65.9733853241, 63.5736445248, 32.944229995, -86.6375999579, 48.3195237109, -54.0662156873, -74.3836623761};
test_label[627] = '{-54.0662156873};
test_output[627] = '{120.126458745};
############ END DEBUG ############*/
test_input[5024:5031] = '{32'h427d85ab, 32'hc282eca3, 32'hc114a57c, 32'hc0db7dd1, 32'h422f34da, 32'h42322a1a, 32'h42554fef, 32'h42a5607d};
test_label[628] = '{32'h42554fef};
test_output[628] = '{32'h41eae215};
/*############ DEBUG ############
test_input[5024:5031] = '{63.3805357652, -65.4621828092, -9.29040128129, -6.85910838016, 43.8016120479, 44.5411139332, 53.328059529, 82.6884512811};
test_label[628] = '{53.328059529};
test_output[628] = '{29.3603917562};
############ END DEBUG ############*/
test_input[5032:5039] = '{32'h42902067, 32'h42ad0d04, 32'h42891992, 32'h3e3fcdc7, 32'h42756feb, 32'hbf3cb51c, 32'hc27b31c5, 32'h41b34394};
test_label[629] = '{32'h42756feb};
test_output[629] = '{32'h41c9543b};
/*############ DEBUG ############
test_input[5032:5039] = '{72.0632868276, 86.5254216095, 68.5499436522, 0.187308420005, 61.3592946453, -0.737138513135, -62.7986012316, 22.407997402};
test_label[629] = '{61.3592946453};
test_output[629] = '{25.1661275037};
############ END DEBUG ############*/
test_input[5040:5047] = '{32'hc272fe6e, 32'h420c0cfe, 32'h42c55b50, 32'h42959684, 32'hc23e13b7, 32'hc0b372b1, 32'h427971fe, 32'hc07c2d44};
test_label[630] = '{32'hc07c2d44};
test_output[630] = '{32'h42cd3cba};
/*############ DEBUG ############
test_input[5040:5047] = '{-60.7484661569, 35.0126891156, 98.678344276, 74.7939723538, -47.5192533649, -5.60775048242, 62.3613202338, -3.94026284788};
test_label[630] = '{-3.94026284788};
test_output[630] = '{102.618607124};
############ END DEBUG ############*/
test_input[5048:5055] = '{32'h4236151f, 32'hc028818e, 32'hc278db19, 32'h415abfaa, 32'h42204ec5, 32'hc270b4d5, 32'hbfccf708, 32'h419b66b7};
test_label[631] = '{32'h415abfaa};
test_output[631] = '{32'h41fed33e};
/*############ DEBUG ############
test_input[5048:5055] = '{45.5206246323, -2.63290744855, -62.2139612578, 13.6717929657, 40.0769239958, -60.1765933643, -1.60128876972, 19.4251539519};
test_label[631] = '{13.6717929657};
test_output[631] = '{31.8531458015};
############ END DEBUG ############*/
test_input[5056:5063] = '{32'hc23b73cf, 32'h42c5af52, 32'hc1c571cc, 32'h4199a3ab, 32'h42b90c02, 32'h42a7a8d0, 32'hc2c3cba3, 32'h42886593};
test_label[632] = '{32'h42c5af52};
test_output[632] = '{32'h3aebfe07};
/*############ DEBUG ############
test_input[5056:5063] = '{-46.8630929485, 98.84242315, -24.6805644344, 19.2049167579, 92.5234530105, 83.8297085328, -97.8977241716, 68.1983843265};
test_label[632] = '{98.84242315};
test_output[632] = '{0.00180047835491};
############ END DEBUG ############*/
test_input[5064:5071] = '{32'hc2c28991, 32'h42986986, 32'hc2078c42, 32'hc21e3ccf, 32'h411f3f5a, 32'hc2686d9d, 32'h4254997b, 32'h4296c088};
test_label[633] = '{32'hc21e3ccf};
test_output[633] = '{32'h42e84135};
/*############ DEBUG ############
test_input[5064:5071] = '{-97.2686873057, 76.2060984783, -33.8869699927, -39.5593826982, 9.95296689162, -58.1070444023, 53.149883099, 75.3760390213};
test_label[633] = '{-39.5593826982};
test_output[633] = '{116.127358915};
############ END DEBUG ############*/
test_input[5072:5079] = '{32'hc1033d00, 32'h4234f3b5, 32'hc2917172, 32'h42463434, 32'hc222f61a, 32'hc288c7d8, 32'hc13e34da, 32'hc20322ac};
test_label[634] = '{32'h42463434};
test_output[634] = '{32'h3c59fb88};
/*############ DEBUG ############
test_input[5072:5079] = '{-8.20239230216, 45.2379935169, -72.7215741936, 49.5509793819, -40.7403317815, -68.3903178358, -11.8879035286, -32.7838610727};
test_label[634] = '{49.5509793819};
test_output[634] = '{0.0133045986566};
############ END DEBUG ############*/
test_input[5080:5087] = '{32'hc256eba0, 32'hc16003a0, 32'hc195e551, 32'h4186e4d4, 32'h41c56c02, 32'hc29b71b4, 32'h42b7f8fa, 32'h42a5d5ba};
test_label[635] = '{32'hc256eba0};
test_output[635] = '{32'h4311b76d};
/*############ DEBUG ############
test_input[5080:5087] = '{-53.7301033934, -14.0008851722, -18.7369713857, 16.8617321529, 24.6777381869, -77.722072953, 91.9862828221, 82.9174360929};
test_label[635] = '{-53.7301033934};
test_output[635] = '{145.716501408};
############ END DEBUG ############*/
test_input[5088:5095] = '{32'hc29ecf4a, 32'hc188318a, 32'hc1f36120, 32'h4097f9b2, 32'hc18092c1, 32'h428baf9a, 32'h42b98379, 32'hc2a5a8f0};
test_label[636] = '{32'hc29ecf4a};
test_output[636] = '{32'h432c2962};
/*############ DEBUG ############
test_input[5088:5095] = '{-79.4048638647, -17.0241882881, -30.4224246629, 4.74923035052, -16.0716581088, 69.8429739267, 92.7567843471, -82.8299527585};
test_label[636] = '{-79.4048638647};
test_output[636] = '{172.161648212};
############ END DEBUG ############*/
test_input[5096:5103] = '{32'h4282fbbe, 32'hc2b5c586, 32'h428ee813, 32'hc28933c3, 32'h40ea8a45, 32'hc29a5633, 32'hc219a708, 32'h42878ea9};
test_label[637] = '{32'hc219a708};
test_output[637] = '{32'h42dbc9b3};
/*############ DEBUG ############
test_input[5096:5103] = '{65.4916868572, -90.8857861968, 71.4532718169, -68.6010991054, 7.32937840376, -77.1683545133, -38.4131174546, 67.7786336076};
test_label[637] = '{-38.4131174546};
test_output[637] = '{109.893940628};
############ END DEBUG ############*/
test_input[5104:5111] = '{32'h42259cc9, 32'hc228828b, 32'hc10cd9de, 32'hc1d9af2f, 32'h424a1fc3, 32'hc299232e, 32'hc20f7834, 32'hc2863fb8};
test_label[638] = '{32'hc2863fb8};
test_output[638] = '{32'h42eb4fa8};
/*############ DEBUG ############
test_input[5104:5111] = '{41.4031086222, -42.1274835522, -8.80319021208, -27.2105396578, 50.5310192046, -76.568709145, -35.8673865114, -67.1244495388};
test_label[638] = '{-67.1244495388};
test_output[638] = '{117.65557733};
############ END DEBUG ############*/
test_input[5112:5119] = '{32'h427243f6, 32'hc2be4b71, 32'h4296fc3b, 32'hc2561e00, 32'hc29a45b6, 32'hc2a79bce, 32'h41099863, 32'hc2ad232b};
test_label[639] = '{32'h41099863};
test_output[639] = '{32'h4285c92f};
/*############ DEBUG ############
test_input[5112:5119] = '{60.5663687721, -95.1473483348, 75.4926401953, -53.5292954968, -77.1361554192, -83.8043042025, 8.59970388, -86.5686875804};
test_label[639] = '{8.59970388};
test_output[639] = '{66.8929366446};
############ END DEBUG ############*/
test_input[5120:5127] = '{32'hc1c67282, 32'h4286f714, 32'hc277f2d1, 32'h42c0ca59, 32'hc1da5f37, 32'h41fb0d38, 32'h42b63776, 32'hc22108e4};
test_label[640] = '{32'hc1c67282};
test_output[640] = '{32'h42f2698f};
/*############ DEBUG ############
test_input[5120:5127] = '{-24.8059120323, 67.4825768899, -61.9871260808, 96.3952113194, -27.2964923202, 31.3814537678, 91.1083244197, -40.2586819286};
test_label[640] = '{-24.8059120323};
test_output[640] = '{121.206168086};
############ END DEBUG ############*/
test_input[5128:5135] = '{32'h41c025a6, 32'hc0f80e7e, 32'h425f5334, 32'h416aa9ef, 32'h3f7d97cc, 32'hbe1058de, 32'hc28d3843, 32'hc20df88a};
test_label[641] = '{32'h425f5334};
test_output[641] = '{32'h288a0000};
/*############ DEBUG ############
test_input[5128:5135] = '{24.0183830341, -7.75176903198, 55.8312520023, 14.6664872801, 0.990597512048, -0.140964006191, -70.6098845184, -35.4927156935};
test_label[641] = '{55.8312520023};
test_output[641] = '{1.53210777398e-14};
############ END DEBUG ############*/
test_input[5136:5143] = '{32'hc2aafe74, 32'hc2c5fe7d, 32'h429cf48a, 32'hc2c35936, 32'h41ec9896, 32'h4220a86c, 32'hc214c8f0, 32'h425bc3e5};
test_label[642] = '{32'hc2c35936};
test_output[642] = '{32'h433026e0};
/*############ DEBUG ############
test_input[5136:5143] = '{-85.4969795954, -98.9970489162, 78.477616241, -97.674240062, 29.5745040592, 40.1644754524, -37.1962297779, 54.9413025886};
test_label[642] = '{-97.674240062};
test_output[642] = '{176.151856303};
############ END DEBUG ############*/
test_input[5144:5151] = '{32'hc2b3f89c, 32'hc2b6b241, 32'h41c1b9f8, 32'hc1d834ed, 32'h428c67ce, 32'h422bb5bf, 32'hc29ec270, 32'hc2c72016};
test_label[643] = '{32'hc2b6b241};
test_output[643] = '{32'h43218d08};
/*############ DEBUG ############
test_input[5144:5151] = '{-89.985563671, -91.3481517741, 24.2158054741, -27.0258419509, 70.2027450536, 42.927484974, -79.3797619682, -99.562664585};
test_label[643] = '{-91.3481517741};
test_output[643] = '{161.550896828};
############ END DEBUG ############*/
test_input[5152:5159] = '{32'h42229eac, 32'h42883c76, 32'h42405af6, 32'h4273099d, 32'h413b1ac7, 32'hc2767e62, 32'hc1e4622f, 32'h425df114};
test_label[644] = '{32'h42405af6};
test_output[644] = '{32'h41a03d3d};
/*############ DEBUG ############
test_input[5152:5159] = '{40.6549517713, 68.118091028, 48.0888290773, 60.7593872959, 11.6940376076, -61.6234205897, -28.5479421513, 55.4854260808};
test_label[644] = '{48.0888290773};
test_output[644] = '{20.0299020352};
############ END DEBUG ############*/
test_input[5160:5167] = '{32'h413f8d93, 32'h42686d79, 32'h41222243, 32'hc28aab6c, 32'h42c46b3d, 32'hc1b9032a, 32'hc2a4e955, 32'hc2b468a3};
test_label[645] = '{32'h413f8d93};
test_output[645] = '{32'h42ac798b};
/*############ DEBUG ############
test_input[5160:5167] = '{11.9720640708, 58.1069065015, 10.1333644015, -69.3348063797, 98.2094513919, -23.1265447609, -82.4557291478, -90.2043652438};
test_label[645] = '{11.9720640708};
test_output[645] = '{86.2373873211};
############ END DEBUG ############*/
test_input[5168:5175] = '{32'hc2a9c50b, 32'h4249379f, 32'h42a4770e, 32'h429be06a, 32'hc11cee0f, 32'h41c81fab, 32'hc112a1ed, 32'hc2948e94};
test_label[646] = '{32'h4249379f};
test_output[646] = '{32'h41ff88bb};
/*############ DEBUG ############
test_input[5168:5175] = '{-84.8848498408, 50.3043172722, 82.2325252376, 77.9383065005, -9.80811994032, 25.015461966, -9.16453281778, -74.2784734703};
test_label[646] = '{50.3043172722};
test_output[646] = '{31.9417629103};
############ END DEBUG ############*/
test_input[5176:5183] = '{32'h42a2cbf5, 32'hc2953bd6, 32'h421c508f, 32'hc28eb8d9, 32'hc2a5afa4, 32'h4125ad1c, 32'hc1b7eeb9, 32'hc259cda6};
test_label[647] = '{32'hc28eb8d9};
test_output[647] = '{32'h4318c267};
/*############ DEBUG ############
test_input[5176:5183] = '{81.3983507436, -74.6168701511, 39.0786712726, -71.3610285311, -82.843049417, 10.3547628096, -22.9915628738, -54.4508268692};
test_label[647] = '{-71.3610285311};
test_output[647] = '{152.759379275};
############ END DEBUG ############*/
test_input[5184:5191] = '{32'hc209bf57, 32'h4191e216, 32'hc22f43fd, 32'h42162f95, 32'h42670bb4, 32'hc0b82822, 32'hc19acd7b, 32'hc2c4affa};
test_label[648] = '{32'hc22f43fd};
test_output[648] = '{32'h42cb27d8};
/*############ DEBUG ############
test_input[5184:5191] = '{-34.4368564923, 18.2353937162, -43.8163950621, 37.5464669668, 57.761427922, -5.75489897303, -19.350332753, -98.3437043808};
test_label[648] = '{-43.8163950621};
test_output[648] = '{101.577822986};
############ END DEBUG ############*/
test_input[5192:5199] = '{32'hc281c1ab, 32'hc2ba2c13, 32'hc299f4d9, 32'h4296ad53, 32'hc251022d, 32'h41bd842e, 32'h41cc48b7, 32'h42a8b8ac};
test_label[649] = '{32'h42a8b8ac};
test_output[649] = '{32'h38fd1ed8};
/*############ DEBUG ############
test_input[5192:5199] = '{-64.8782585176, -93.086083061, -76.9782203308, 75.3385237706, -52.2521265819, 23.6895403347, 25.5355053654, 84.3606885978};
test_label[649] = '{84.3606885978};
test_output[649] = '{0.000120697254514};
############ END DEBUG ############*/
test_input[5200:5207] = '{32'h42c18ee3, 32'hc2b395e7, 32'h42ab0204, 32'hc1245875, 32'h42920d53, 32'h42824e70, 32'hc27b8578, 32'h4152ac9a};
test_label[650] = '{32'h42c18ee3};
test_output[650] = '{32'h3754ceed};
/*############ DEBUG ############
test_input[5200:5207] = '{96.7790745316, -89.7927810069, 85.5039364805, -10.2715961763, 73.0260204545, 65.1531975162, -62.8803396199, 13.1671391956};
test_label[650] = '{96.7790745316};
test_output[650] = '{1.26843630118e-05};
############ END DEBUG ############*/
test_input[5208:5215] = '{32'hc09388c0, 32'hc29b03f2, 32'h42876700, 32'h410edf0f, 32'h400b8ad1, 32'hc2285a07, 32'h4297036e, 32'h42bf80f2};
test_label[651] = '{32'h42bf80f2};
test_output[651] = '{32'h30ddc89a};
/*############ DEBUG ############
test_input[5208:5215] = '{-4.61044326175, -77.5077075503, 67.7011732553, 8.92945801637, 2.18034761769, -42.0879160482, 75.5066977918, 95.7518486773};
test_label[651] = '{95.7518486773};
test_output[651] = '{1.61368807336e-09};
############ END DEBUG ############*/
test_input[5216:5223] = '{32'h4142b89d, 32'hc2acbdae, 32'hc1a537d4, 32'hc1c7c613, 32'h42847026, 32'hc238db47, 32'hc25f0781, 32'h4274c056};
test_label[652] = '{32'hc238db47};
test_output[652] = '{32'h42e0e11f};
/*############ DEBUG ############
test_input[5216:5223] = '{12.1700714166, -86.3704684951, -20.652259096, -24.9717165977, 66.2190432351, -46.2141382958, -55.7573261599, 61.1878274734};
test_label[652] = '{-46.2141382958};
test_output[652] = '{112.439691163};
############ END DEBUG ############*/
test_input[5224:5231] = '{32'hc28c1165, 32'h4287dec9, 32'h4292463b, 32'hc0b8c6f0, 32'hc1a54bd5, 32'hc2b4b489, 32'h422fe888, 32'hc1bfeb1f};
test_label[653] = '{32'hc0b8c6f0};
test_output[653] = '{32'h429dd57a};
/*############ DEBUG ############
test_input[5224:5231] = '{-70.0339744436, 67.935124395, 73.137172489, -5.77428451935, -20.6620267512, -90.3526063284, 43.9770821721, -23.989805921};
test_label[653] = '{-5.77428451935};
test_output[653] = '{78.9169471873};
############ END DEBUG ############*/
test_input[5232:5239] = '{32'hc1b58a85, 32'h4190580a, 32'hc21dd01c, 32'hc2a11925, 32'h426efddf, 32'hc2c62099, 32'hc24a38a0, 32'h4235db7d};
test_label[654] = '{32'hc1b58a85};
test_output[654] = '{32'h42a4e191};
/*############ DEBUG ############
test_input[5232:5239] = '{-22.6926371806, 18.0429876034, -39.4532300591, -80.5491135704, 59.7479221491, -99.0636689059, -50.5552996988, 45.4643441688};
test_label[654] = '{-22.6926371806};
test_output[654] = '{82.4405599559};
############ END DEBUG ############*/
test_input[5240:5247] = '{32'hbf06a025, 32'hc26bb37d, 32'hc252490b, 32'hc206476e, 32'hc220c7b1, 32'h422cfa6c, 32'hc2443ae9, 32'hc1181bb1};
test_label[655] = '{32'hc26bb37d};
test_output[655] = '{32'h42cc56f5};
/*############ DEBUG ############
test_input[5240:5247] = '{-0.525881127228, -58.9252826495, -52.5713291504, -33.5697552379, -40.1950115997, 43.2445543775, -49.0575285921, -9.50676068176};
test_label[655] = '{-58.9252826495};
test_output[655] = '{102.169837027};
############ END DEBUG ############*/
test_input[5248:5255] = '{32'hc1947ef3, 32'hc0ea7499, 32'h41994117, 32'h41851b8b, 32'hc2497596, 32'hc2055cd3, 32'h4218937e, 32'hc1f26152};
test_label[656] = '{32'hc0ea7499};
test_output[656] = '{32'h4235e211};
/*############ DEBUG ############
test_input[5248:5255] = '{-18.5619869116, -7.32673316804, 19.156781543, 16.6384488939, -50.3648284501, -33.3406493708, 38.1440339517, -30.2975204413};
test_label[656] = '{-7.32673316804};
test_output[656] = '{45.4707671259};
############ END DEBUG ############*/
test_input[5256:5263] = '{32'hc265fe76, 32'h42669c97, 32'hc1a53bd0, 32'hc2984977, 32'hc05fd023, 32'hc2b5669e, 32'hc2961e49, 32'h42868fcf};
test_label[657] = '{32'h42868fcf};
test_output[657] = '{32'h388a1df5};
/*############ DEBUG ############
test_input[5256:5263] = '{-57.498495373, 57.6529182316, -20.6542045742, -76.1434870277, -3.49707872169, -90.7004271391, -75.0591512231, 67.2808748108};
test_label[657] = '{67.2808748108};
test_output[657] = '{6.5859326383e-05};
############ END DEBUG ############*/
test_input[5264:5271] = '{32'hc0d04bd1, 32'h41d3ddb9, 32'hc20edaa5, 32'hc26c17f5, 32'hc1d2eda1, 32'hc1dbf406, 32'hc20b7282, 32'h41b17a55};
test_label[658] = '{32'h41d3ddb9};
test_output[658] = '{32'h3c5d229d};
/*############ DEBUG ############
test_input[5264:5271] = '{-6.50925497392, 26.4832626551, -35.7135196166, -59.0233936887, -26.3660291669, -27.4941528087, -34.861822445, 22.1847325119};
test_label[658] = '{26.4832626551};
test_output[658] = '{0.0134970215421};
############ END DEBUG ############*/
test_input[5272:5279] = '{32'h41eb5ab3, 32'h421e3a0b, 32'h42388e22, 32'h429f56c0, 32'h42a81cf5, 32'hc1db654e, 32'hc186b383, 32'hc200bb9c};
test_label[659] = '{32'h421e3a0b};
test_output[659] = '{32'h42320c86};
/*############ DEBUG ############
test_input[5272:5279] = '{29.4192865993, 39.5566833986, 46.1388011122, 79.6694343569, 84.0565535779, -27.4244645973, -16.8376515513, -32.1832112678};
test_label[659] = '{39.5566833986};
test_output[659] = '{44.5122299857};
############ END DEBUG ############*/
test_input[5280:5287] = '{32'hc291dc8a, 32'hc22474d5, 32'hc1ac66b2, 32'h41e627da, 32'hc1ef4cf4, 32'h4296e28d, 32'h41f88c41, 32'hc235eeb5};
test_label[660] = '{32'h4296e28d};
test_output[660] = '{32'h80000000};
/*############ DEBUG ############
test_input[5280:5287] = '{-72.9307400221, -41.1140941589, -21.5501434193, 28.7694582449, -29.912573964, 75.4424815849, 31.0684826223, -45.4831108474};
test_label[660] = '{75.4424815849};
test_output[660] = '{-0.0};
############ END DEBUG ############*/
test_input[5288:5295] = '{32'h428e1db3, 32'hc195b116, 32'h402ad323, 32'h41f58164, 32'h415f5c35, 32'h42358c72, 32'hc2b05756, 32'h42adca90};
test_label[661] = '{32'h415f5c35};
test_output[661] = '{32'h4291df0a};
/*############ DEBUG ############
test_input[5288:5295] = '{71.0580031154, -18.7114675073, 2.66913667959, 30.6881798029, 13.9600117136, 45.3871528988, -88.1705804603, 86.8956317763};
test_label[661] = '{13.9600117136};
test_output[661] = '{72.935620195};
############ END DEBUG ############*/
test_input[5296:5303] = '{32'hc179e8cd, 32'hc0a2984d, 32'hc161f6c1, 32'hc2ba8d62, 32'h41759dbe, 32'hc2aaf52b, 32'hc184bcf4, 32'hc201e72f};
test_label[662] = '{32'h41759dbe};
test_output[662] = '{32'h30b7eb63};
/*############ DEBUG ############
test_input[5296:5303] = '{-15.6193363599, -5.08109164205, -14.1227425765, -93.2761391105, 15.3510108198, -85.4788474055, -16.5922621857, -32.4757665837};
test_label[662] = '{15.3510108198};
test_output[662] = '{1.33819033722e-09};
############ END DEBUG ############*/
test_input[5304:5311] = '{32'h42bfbd2c, 32'hc27a2a05, 32'hc194cdf8, 32'h40cecaef, 32'hc2133550, 32'hc24fe0aa, 32'hc2753f0b, 32'h41b2a006};
test_label[663] = '{32'hc27a2a05};
test_output[663] = '{32'h431e6918};
/*############ DEBUG ############
test_input[5304:5311] = '{95.8694792638, -62.541035989, -18.6005699429, 6.46227229718, -36.8020626188, -51.9693988079, -61.3115637921, 22.3281366118};
test_label[663] = '{-62.541035989};
test_output[663] = '{158.410515253};
############ END DEBUG ############*/
test_input[5312:5319] = '{32'hc2c33a99, 32'hc141e270, 32'h428c1855, 32'h40089f5a, 32'h423ca6f1, 32'h40b2ca14, 32'hc299c468, 32'hc299867b};
test_label[664] = '{32'hc2c33a99};
test_output[664] = '{32'h4327a977};
/*############ DEBUG ############
test_input[5312:5319] = '{-97.6144459581, -12.1177823105, 70.0475215868, 2.13472607646, 47.163027575, 5.58716771344, -76.8836054047, -76.7626572183};
test_label[664] = '{-97.6144459581};
test_output[664] = '{167.661967545};
############ END DEBUG ############*/
test_input[5320:5327] = '{32'h400b6cba, 32'h429e6457, 32'h42a86b9e, 32'h419420ea, 32'h42993b9c, 32'h40d056ae, 32'hc1c486e4, 32'h428e7db1};
test_label[665] = '{32'h42a86b9e};
test_output[665] = '{32'h3be96aec};
/*############ DEBUG ############
test_input[5320:5327] = '{2.17851110656, 79.1959751685, 84.2101892117, 18.5160713114, 76.6164222546, 6.51058092671, -24.5658642835, 71.2454902743};
test_label[665] = '{84.2101892117};
test_output[665] = '{0.0071233416892};
############ END DEBUG ############*/
test_input[5328:5335] = '{32'hc2b37c84, 32'hc27fa899, 32'h40a55ec3, 32'h41102cdd, 32'hc1b1fe29, 32'hc24d9c25, 32'h415b7b32, 32'h423e1aac};
test_label[666] = '{32'h40a55ec3};
test_output[666] = '{32'h42296ed4};
/*############ DEBUG ############
test_input[5328:5335] = '{-89.7431961751, -63.9146446189, 5.16781748839, 9.01095247723, -22.2491021616, -51.402484415, 13.7175767384, 47.5260461968};
test_label[666] = '{5.16781748839};
test_output[666] = '{42.3582287085};
############ END DEBUG ############*/
test_input[5336:5343] = '{32'h4189bbc8, 32'h41c4036b, 32'hc26c7877, 32'hc276f29a, 32'h42979fc1, 32'hc2839c21, 32'h418ef43c, 32'h3fcd53a0};
test_label[667] = '{32'h42979fc1};
test_output[667] = '{32'h80000000};
/*############ DEBUG ############
test_input[5336:5343] = '{17.2166907603, 24.501668613, -59.1176404308, -61.7369147948, 75.8120165463, -65.8049393207, 17.869255388, 1.60411451459};
test_label[667] = '{75.8120165463};
test_output[667] = '{-0.0};
############ END DEBUG ############*/
test_input[5344:5351] = '{32'hc1022b94, 32'h42a69e2c, 32'hc24e0f26, 32'h42ae0b31, 32'h427b773f, 32'h400890ff, 32'h41ea7df7, 32'h42aaaeeb};
test_label[668] = '{32'h427b773f};
test_output[668] = '{32'h41c2c5ea};
/*############ DEBUG ############
test_input[5344:5351] = '{-8.13563900959, 83.3089308747, -51.5147947997, 87.0218586102, 62.8664519706, 2.1338499354, 29.311506047, 85.341640196};
test_label[668] = '{62.8664519706};
test_output[668] = '{24.3466377532};
############ END DEBUG ############*/
test_input[5352:5359] = '{32'h40e74907, 32'h40dbe7f1, 32'h426b338c, 32'h41d7ed21, 32'h42045dec, 32'hc25c5861, 32'hc205f3ff, 32'h4112e35d};
test_label[669] = '{32'hc25c5861};
test_output[669] = '{32'h42e3c5f6};
/*############ DEBUG ############
test_input[5352:5359] = '{7.22766465742, 6.87206336515, 58.8003400146, 26.9907862355, 33.0917191064, -55.0863061664, -33.4882761014, 9.18050826444};
test_label[669] = '{-55.0863061664};
test_output[669] = '{113.886646181};
############ END DEBUG ############*/
test_input[5360:5367] = '{32'hc1855af0, 32'hc2bcdc92, 32'hc29cf4ba, 32'h41d3b909, 32'h41a1dceb, 32'h423410ee, 32'h412dfb07, 32'hc1df7cb4};
test_label[670] = '{32'hc1855af0};
test_output[670] = '{32'h4276be66};
/*############ DEBUG ############
test_input[5360:5367] = '{-16.6694027796, -94.430799263, -78.4779789933, 26.4653484974, 20.2328703472, 45.0165346725, 10.8737858649, -27.9358899368};
test_label[670] = '{-16.6694027796};
test_output[670] = '{61.6859374609};
############ END DEBUG ############*/
test_input[5368:5375] = '{32'h40d09337, 32'hc2412e45, 32'hc2a217d4, 32'h4287c691, 32'hc20235f5, 32'h4232e150, 32'h4236fa8e, 32'h41cc4abd};
test_label[671] = '{32'h40d09337};
test_output[671] = '{32'h42757abb};
/*############ DEBUG ############
test_input[5368:5375] = '{6.51797062008, -48.2951847948, -81.046536636, 67.8878246999, -32.552691286, 44.7200332117, 45.7446833842, 25.536493801};
test_label[671] = '{6.51797062008};
test_output[671] = '{61.3698540801};
############ END DEBUG ############*/
test_input[5376:5383] = '{32'h410362a0, 32'h42b2471e, 32'h42add131, 32'h41836f0c, 32'hc14bd94c, 32'hc0e36120, 32'h42290ab8, 32'h42388759};
test_label[672] = '{32'hc14bd94c};
test_output[672] = '{32'h42cbf68e};
/*############ DEBUG ############
test_input[5376:5383] = '{8.21157807659, 89.1389021332, 86.908580242, 16.4292214637, -12.7405512784, -7.10560622217, 42.2604658235, 46.1321738684};
test_label[672] = '{-12.7405512784};
test_output[672] = '{101.981553057};
############ END DEBUG ############*/
test_input[5384:5391] = '{32'h4290872e, 32'h42acb2c0, 32'h429cd1df, 32'h4255f50e, 32'h428356cf, 32'hbf1a99e3, 32'hc296f79b, 32'hc1645315};
test_label[673] = '{32'h429cd1df};
test_output[673] = '{32'h40fe1100};
/*############ DEBUG ############
test_input[5384:5391] = '{72.2640210097, 86.3491227132, 78.4099048213, 53.4893123413, 65.669551817, -0.603910639013, -75.483607553, -14.2702841076};
test_label[673] = '{78.4099048213};
test_output[673] = '{7.93957507802};
############ END DEBUG ############*/
test_input[5392:5399] = '{32'hc2b61cfa, 32'hc23cc0b0, 32'h41adbe73, 32'h41293637, 32'h429b9cb8, 32'hc2658740, 32'h4236cdb3, 32'hc2afb7e8};
test_label[674] = '{32'h41adbe73};
test_output[674] = '{32'h42605a37};
/*############ DEBUG ############
test_input[5392:5399] = '{-91.0565949064, -47.1881723102, 21.7179930852, 10.5757359596, 77.8060947462, -57.3820795647, 45.7008774838, -87.8591893845};
test_label[674] = '{21.7179930852};
test_output[674] = '{56.088101661};
############ END DEBUG ############*/
test_input[5400:5407] = '{32'hc129a990, 32'h41c01758, 32'h42a8117a, 32'hc25bcd38, 32'hc2822225, 32'h42ae50f3, 32'h41c44337, 32'h42712011};
test_label[675] = '{32'h42ae50f3};
test_output[675] = '{32'h3d304d60};
/*############ DEBUG ############
test_input[5400:5407] = '{-10.6038971819, 24.0113984375, 84.034135507, -54.9504084063, -65.0666920113, 87.1581034123, 24.532819316, 60.2813144313};
test_label[675] = '{87.1581034123};
test_output[675] = '{0.0430425392335};
############ END DEBUG ############*/
test_input[5408:5415] = '{32'h42bfcc5d, 32'h420deaf0, 32'h42c47aa3, 32'h42938db3, 32'h42a1b374, 32'h42815b1c, 32'hc23380eb, 32'hc1638778};
test_label[676] = '{32'h42a1b374};
test_output[676] = '{32'h418bd903};
/*############ DEBUG ############
test_input[5408:5415] = '{95.8991483088, 35.4794300666, 98.2395217866, 73.7767570771, 80.850493056, 64.6779493003, -44.875895129, -14.2205732151};
test_label[676] = '{80.850493056};
test_output[676] = '{17.4809620304};
############ END DEBUG ############*/
test_input[5416:5423] = '{32'hc2af936c, 32'hc1f49ec6, 32'h416668a4, 32'h4216eaca, 32'h42bf3fd8, 32'h427fefc2, 32'hc10750bf, 32'hc16f910a};
test_label[677] = '{32'h42bf3fd8};
test_output[677] = '{32'h28a40000};
/*############ DEBUG ############
test_input[5416:5423] = '{-87.7879325228, -30.5775257598, 14.4005467505, 37.7292847711, 95.6246918329, 63.9841387456, -8.45721322043, -14.9729103121};
test_label[677] = '{95.6246918329};
test_output[677] = '{1.82076576039e-14};
############ END DEBUG ############*/
test_input[5424:5431] = '{32'hc17a1d16, 32'hc26c9088, 32'hc1f49278, 32'h426cd915, 32'h42b9fe9f, 32'h41cb7e57, 32'hc1e9e9d9, 32'hc244a587};
test_label[678] = '{32'hc26c9088};
test_output[678] = '{32'h43182372};
/*############ DEBUG ############
test_input[5424:5431] = '{-15.6321009273, -59.1411424521, -30.5715184958, 59.2119959092, 92.9973090932, 25.4366902571, -29.2391840067, -49.1616482327};
test_label[678] = '{-59.1411424521};
test_output[678] = '{152.138451545};
############ END DEBUG ############*/
test_input[5432:5439] = '{32'h423a632a, 32'h42abc107, 32'h42bd9970, 32'hc2b8122e, 32'hbfd49fac, 32'hc1dac83f, 32'hc28d94bb, 32'h42a0853c};
test_label[679] = '{32'h42a0853c};
test_output[679] = '{32'h4168a22b};
/*############ DEBUG ############
test_input[5432:5439] = '{46.5968407616, 85.8770082574, 94.7996824405, -92.0355102912, -1.66112285347, -27.3477773176, -70.790486765, 80.2602243391};
test_label[679] = '{80.2602243391};
test_output[679] = '{14.5395919086};
############ END DEBUG ############*/
test_input[5440:5447] = '{32'hc24c5c34, 32'hc2b3ba7e, 32'h42aed968, 32'h4286ede7, 32'hc23bfca5, 32'h42a56615, 32'hc123becd, 32'hc1316ec0};
test_label[680] = '{32'h42a56615};
test_output[680] = '{32'h40977d7c};
/*############ DEBUG ############
test_input[5440:5447] = '{-51.0900416062, -89.8642462882, 87.4246197027, 67.4646539171, -46.9967228924, 82.6993813932, -10.2340826855, -11.0895387144};
test_label[680] = '{82.6993813932};
test_output[680] = '{4.73406781681};
############ END DEBUG ############*/
test_input[5448:5455] = '{32'h424229e4, 32'h429c621a, 32'hc0b42402, 32'h4206aa45, 32'hc00b9316, 32'h4183d00a, 32'h40b0271a, 32'h42a6681f};
test_label[681] = '{32'h4183d00a};
test_output[681] = '{32'h42857783};
/*############ DEBUG ############
test_input[5448:5455] = '{48.5409100177, 78.1916015893, -5.62939546753, 33.6662787911, -2.18085252224, 16.4765819645, 5.50477301803, 83.2033638313};
test_label[681] = '{16.4765819645};
test_output[681] = '{66.7334189504};
############ END DEBUG ############*/
test_input[5456:5463] = '{32'hc238d187, 32'h426e62a5, 32'hc269d3e7, 32'h40a5e0fe, 32'h4281a0bb, 32'h417ba2c5, 32'h42329f9c, 32'h429da98c};
test_label[682] = '{32'hc238d187};
test_output[682] = '{32'h42fa1250};
/*############ DEBUG ############
test_input[5456:5463] = '{-46.2046149204, 59.5963313183, -58.4569375223, 5.18371466367, 64.8139276996, 15.7272390721, 44.6558677132, 78.8311492414};
test_label[682] = '{-46.2046149204};
test_output[682] = '{125.035764984};
############ END DEBUG ############*/
test_input[5464:5471] = '{32'hc2b6f774, 32'h421d3dd7, 32'h422d08a8, 32'hc2abf647, 32'hc1d3ea9c, 32'h42963ae8, 32'h422f1f4c, 32'hc1b192f2};
test_label[683] = '{32'hc2b6f774};
test_output[683] = '{32'h4326992e};
/*############ DEBUG ############
test_input[5464:5471] = '{-91.4833101279, 39.3103896475, 43.2584532592, -85.9810079287, -26.4895558962, 75.1150498074, 43.7805642648, -22.1967508054};
test_label[683] = '{-91.4833101279};
test_output[683] = '{166.598359935};
############ END DEBUG ############*/
test_input[5472:5479] = '{32'hc2b0b704, 32'hc2a60c15, 32'h429a7cc7, 32'h42aae206, 32'h42a5f187, 32'hc2545eef, 32'hc2170d60, 32'h41adf2e1};
test_label[684] = '{32'h41adf2e1};
test_output[684] = '{32'h427f1e09};
/*############ DEBUG ############
test_input[5472:5479] = '{-88.3574561412, -83.023594954, 77.2437083221, 85.441450794, 82.9717340857, -53.0927091649, -37.7630628969, 21.7435924214};
test_label[684] = '{21.7435924214};
test_output[684] = '{63.7793315326};
############ END DEBUG ############*/
test_input[5480:5487] = '{32'h41b3405f, 32'hc2c64a6e, 32'hc2005fa9, 32'h41d59eb6, 32'hc2acf502, 32'h4077963f, 32'h415036d4, 32'h4093f20f};
test_label[685] = '{32'h415036d4};
test_output[685] = '{32'h415b3e05};
/*############ DEBUG ############
test_input[5480:5487] = '{22.4064318858, -99.1453740304, -32.0934185905, 26.7024956653, -86.4785301784, 3.86854540782, 13.0133854175, 4.62329798594};
test_label[685] = '{13.0133854175};
test_output[685] = '{13.7026414945};
############ END DEBUG ############*/
test_input[5488:5495] = '{32'hc25e69cb, 32'h42590f9a, 32'h428fc9fc, 32'h42b4cbb0, 32'hc1f7b53b, 32'hc270c7fa, 32'hc17059b2, 32'h42c6aab5};
test_label[686] = '{32'hc1f7b53b};
test_output[686] = '{32'h43024c0a};
/*############ DEBUG ############
test_input[5488:5495] = '{-55.6033119697, 54.2652346262, 71.8945004483, 90.3978252697, -30.9634923865, -60.1952906863, -15.0218979242, 99.3334085843};
test_label[686] = '{-30.9634923865};
test_output[686] = '{130.297032583};
############ END DEBUG ############*/
test_input[5496:5503] = '{32'h41c178c1, 32'hc2b0752a, 32'h42263b8b, 32'h42015678, 32'hc1ede094, 32'h429e224c, 32'h41409b46, 32'h41ee74b2};
test_label[687] = '{32'h41ee74b2};
test_output[687] = '{32'h42450a3f};
/*############ DEBUG ############
test_input[5496:5503] = '{24.1839627285, -88.2288323432, 41.5581476817, 32.3344436005, -29.7346569051, 79.0669868533, 12.0379087832, 29.8069800687};
test_label[687] = '{29.8069800687};
test_output[687] = '{49.2600067847};
############ END DEBUG ############*/
test_input[5504:5511] = '{32'hc289805c, 32'hc24653ce, 32'hc19b4393, 32'hc2078e25, 32'h425f4f7d, 32'h42b68f63, 32'h42483579, 32'hc28b9595};
test_label[688] = '{32'hc2078e25};
test_output[688] = '{32'h42fa5676};
/*############ DEBUG ############
test_input[5504:5511] = '{-68.7507054149, -49.5818394118, -19.4079950375, -33.888814703, 55.8276260485, 91.280050679, 50.0522191835, -69.7921489667};
test_label[688] = '{-33.888814703};
test_output[688] = '{125.168865382};
############ END DEBUG ############*/
test_input[5512:5519] = '{32'hc1acc189, 32'hc2c6a8d5, 32'hc29f244d, 32'h42b7c34c, 32'h40b7276c, 32'hc2394929, 32'hc2aa5bb9, 32'h420c470f};
test_label[689] = '{32'h420c470f};
test_output[689] = '{32'h42633f8a};
/*############ DEBUG ############
test_input[5512:5519] = '{-21.5945002837, -99.3297524956, -79.5709007198, 91.8814423384, 5.72356225449, -46.321444925, -85.1791421365, 35.0693914468};
test_label[689] = '{35.0693914468};
test_output[689] = '{56.8120508916};
############ END DEBUG ############*/
test_input[5520:5527] = '{32'hc2854e16, 32'hc29cd8a5, 32'h4245ce7c, 32'hc2ba3dff, 32'hc2815c93, 32'hc259f3d9, 32'h4010bedd, 32'hc25507fa};
test_label[690] = '{32'hc259f3d9};
test_output[690] = '{32'h42cfe12b};
/*############ DEBUG ############
test_input[5520:5527] = '{-66.6525139771, -78.4231323689, 49.4516448006, -93.1210887359, -64.6808088921, -54.4881327736, 2.26164944129, -53.2577913409};
test_label[690] = '{-54.4881327736};
test_output[690] = '{103.939777574};
############ END DEBUG ############*/
test_input[5528:5535] = '{32'hc28aadf4, 32'hc2543fda, 32'h42c78a87, 32'h429961b3, 32'h41928f6c, 32'hc1931ff8, 32'h42852add, 32'hc280790a};
test_label[691] = '{32'h42852add};
test_output[691] = '{32'h4204bf55};
/*############ DEBUG ############
test_input[5528:5535] = '{-69.3397523875, -53.0623561876, 99.7705643565, 76.6908207968, 18.3200294816, -18.3906095305, 66.5837175751, -64.2364060676};
test_label[691] = '{66.5837175751};
test_output[691] = '{33.1868467815};
############ END DEBUG ############*/
test_input[5536:5543] = '{32'h419402c9, 32'h428b9c14, 32'hc23e06b4, 32'h42c48435, 32'h42874bd2, 32'h4208b2fd, 32'hc181709f, 32'h428057df};
test_label[692] = '{32'h42c48435};
test_output[692] = '{32'h2b0a7000};
/*############ DEBUG ############
test_input[5536:5543] = '{18.5013605258, 69.8048383756, -47.5065467318, 98.2582151035, 67.6480877898, 34.1747927901, -16.1799903068, 64.1716240704};
test_label[692] = '{98.2582151035};
test_output[692] = '{4.91828799909e-13};
############ END DEBUG ############*/
test_input[5544:5551] = '{32'h428ffa26, 32'h403e64ef, 32'hc216c1ff, 32'hc2a36878, 32'hc202e18d, 32'h420a74ae, 32'h4226b407, 32'hc20f62e4};
test_label[693] = '{32'h428ffa26};
test_output[693] = '{32'h299a4000};
/*############ DEBUG ############
test_input[5544:5551] = '{71.9885725141, 2.97491056387, -37.6894487803, -81.7040416847, -32.7202646166, 34.6139437491, 41.6758098478, -35.8465734308};
test_label[693] = '{71.9885725141};
test_output[693] = '{6.85007606194e-14};
############ END DEBUG ############*/
test_input[5552:5559] = '{32'h41c7b425, 32'h4246f77d, 32'h42bf36cb, 32'h428df934, 32'hc286e848, 32'h428318a7, 32'h42a0d2f9, 32'hc1b5980e};
test_label[694] = '{32'h42a0d2f9};
test_output[694] = '{32'h41731e91};
/*############ DEBUG ############
test_input[5552:5559] = '{24.9629611619, 49.7416871146, 95.6070205129, 70.9867267554, -67.45367772, 65.5481481701, 80.4120583176, -22.6992459009};
test_label[694] = '{80.4120583176};
test_output[694] = '{15.194962447};
############ END DEBUG ############*/
test_input[5560:5567] = '{32'h40a68590, 32'hc2ab5ef8, 32'hc23ea143, 32'h4275aead, 32'hc2911be6, 32'h42aee25c, 32'hc23815a0, 32'h40a27522};
test_label[695] = '{32'h4275aead};
test_output[695] = '{32'h41d02c15};
/*############ DEBUG ############
test_input[5560:5567] = '{5.20380411543, -85.6854869767, -47.6574828704, 61.4205834452, -72.5544888093, 87.4421077667, -46.0211195439, 5.07679854813};
test_label[695] = '{61.4205834452};
test_output[695] = '{26.0215243215};
############ END DEBUG ############*/
test_input[5568:5575] = '{32'hc2aa4401, 32'h40beef06, 32'hc2bf0e6d, 32'hc29a87cd, 32'hc1b1426c, 32'h42118349, 32'h4246dff6, 32'hc18e94f9};
test_label[696] = '{32'h4246dff6};
test_output[696] = '{32'h35d7d35d};
/*############ DEBUG ############
test_input[5568:5575] = '{-85.1328205077, 5.96667754954, -95.528178748, -77.2652339357, -22.1574333882, 36.3782079251, 49.7187101137, -17.8227414313};
test_label[696] = '{49.7187101137};
test_output[696] = '{1.60802636286e-06};
############ END DEBUG ############*/
test_input[5576:5583] = '{32'h41ae33c8, 32'hc2815e52, 32'hc1676b27, 32'hc29bc424, 32'hc2776e4f, 32'hc21e5ea0, 32'hc1db7bdf, 32'hc285aa5a};
test_label[697] = '{32'hc285aa5a};
test_output[697] = '{32'h42b1374b};
/*############ DEBUG ############
test_input[5576:5583] = '{21.7752828746, -64.6842173696, -14.4636605508, -77.8830846754, -61.8577246997, -39.5924062374, -27.4354842293, -66.8327141588};
test_label[697] = '{-66.8327141588};
test_output[697] = '{88.6079970334};
############ END DEBUG ############*/
test_input[5584:5591] = '{32'hc2715a2c, 32'h427f2789, 32'h42b5b0f2, 32'hc2c63761, 32'h41d24072, 32'hc29f46ee, 32'hc1e08dfd, 32'h42092a5e};
test_label[698] = '{32'hc29f46ee};
test_output[698] = '{32'h432a7bf0};
/*############ DEBUG ############
test_input[5584:5591] = '{-60.3380593795, 63.7886093558, 90.8455939666, -99.1081606715, 26.2814675996, -79.6385362919, -28.0693299639, 34.2913729834};
test_label[698] = '{-79.6385362919};
test_output[698] = '{170.484130258};
############ END DEBUG ############*/
test_input[5592:5599] = '{32'h40a1bfd9, 32'h413bf8d1, 32'h429f5d3b, 32'hc2226902, 32'hc2be07cb, 32'h4289ce37, 32'h42bf0ba8, 32'h42c182fe};
test_label[699] = '{32'hc2be07cb};
test_output[699] = '{32'h434006dc};
/*############ DEBUG ############
test_input[5592:5599] = '{5.05466880441, 11.7482457749, 79.6820943523, -40.602547441, -95.015224119, 68.9027625973, 95.5227625995, 96.7558407183};
test_label[699] = '{-95.015224119};
test_output[699] = '{192.026787315};
############ END DEBUG ############*/
test_input[5600:5607] = '{32'hc220be6d, 32'h42976382, 32'hc1bc289b, 32'hbf2c5ff5, 32'h42b53fe8, 32'hc2b11d78, 32'h41ef42c2, 32'hc28ea7cf};
test_label[700] = '{32'h42b53fe8};
test_output[700] = '{32'h34b00e8a};
/*############ DEBUG ############
test_input[5600:5607] = '{-40.185962297, 75.6943519358, -23.5198266391, -0.673339159983, 90.6248133972, -88.5575536412, 29.907597153, -71.3277517555};
test_label[700] = '{90.6248133972};
test_output[700] = '{3.27931325018e-07};
############ END DEBUG ############*/
test_input[5608:5615] = '{32'hc111b45a, 32'hc29119d6, 32'hc1f532d0, 32'hc1e00a07, 32'h412b2774, 32'hc263a94b, 32'hc281fa40, 32'h4048f68f};
test_label[701] = '{32'hc29119d6};
test_output[701] = '{32'h42a67f09};
/*############ DEBUG ############
test_input[5608:5615] = '{-9.10653159793, -72.5504621187, -30.6498106518, -28.0048960978, 10.6971320158, -56.9153252813, -64.9887702709, 3.14004883049};
test_label[701] = '{-72.5504621187};
test_output[701] = '{83.2481163974};
############ END DEBUG ############*/
test_input[5616:5623] = '{32'h42882f46, 32'hc2bc09f1, 32'hc2af6d88, 32'h423dd352, 32'hc20741fe, 32'h42704da2, 32'h4223f061, 32'h42bc48e1};
test_label[702] = '{32'h42882f46};
test_output[702] = '{32'h41d0666a};
/*############ DEBUG ############
test_input[5616:5623] = '{68.092332427, -94.0194132286, -87.7139258321, 47.4563690797, -33.814445588, 60.0758141048, 40.9847437775, 94.1423401274};
test_label[702] = '{68.092332427};
test_output[702] = '{26.0500077005};
############ END DEBUG ############*/
test_input[5624:5631] = '{32'hc0d59b4b, 32'h42ac6fbc, 32'hc28c9fed, 32'h42b2b878, 32'h42967268, 32'h41a50c00, 32'h42063897, 32'h4196fb74};
test_label[703] = '{32'h41a50c00};
test_output[703] = '{32'h42898b1e};
/*############ DEBUG ############
test_input[5624:5631] = '{-6.67520685996, 86.2182333286, -70.3123536935, 89.3602872388, 75.2234474219, 20.6308594467, 33.555264692, 18.8727799218};
test_label[703] = '{20.6308594467};
test_output[703] = '{68.7717156384};
############ END DEBUG ############*/
test_input[5632:5639] = '{32'hc29a255c, 32'h420e6b14, 32'hc180b062, 32'h41ab11b1, 32'h42b92585, 32'hc2a8b08d, 32'hc2b347fc, 32'hc2118079};
test_label[704] = '{32'hc29a255c};
test_output[704] = '{32'h4329a571};
/*############ DEBUG ############
test_input[5632:5639] = '{-77.0729690643, 35.6045700293, -16.086125295, 21.3836378062, 92.5732825704, -84.3448235297, -89.6405938302, -36.3754604836};
test_label[704] = '{-77.0729690643};
test_output[704] = '{169.646251635};
############ END DEBUG ############*/
test_input[5640:5647] = '{32'hc2af8b29, 32'hc26eacd1, 32'hbed3d0cd, 32'h41bdc533, 32'hc118be03, 32'h42251f67, 32'h42c08ae9, 32'hc1f3ce46};
test_label[705] = '{32'hc26eacd1};
test_output[705] = '{32'h431bf0a9};
/*############ DEBUG ############
test_input[5640:5647] = '{-87.7717958458, -59.6687648785, -0.413702409188, 23.7212882784, -9.5463899957, 41.2806672851, 96.2713110544, -30.4757189968};
test_label[705] = '{-59.6687648785};
test_output[705] = '{155.940075933};
############ END DEBUG ############*/
test_input[5648:5655] = '{32'hc08075d6, 32'hc1c54cd0, 32'hc11be6ac, 32'hc1bf0da1, 32'h42649965, 32'hc1bac27e, 32'hc2c32af5, 32'hc272f09f};
test_label[706] = '{32'hc08075d6};
test_output[706] = '{32'h4274a81f};
/*############ DEBUG ############
test_input[5648:5655] = '{-4.0143842342, -24.6625064236, -9.74381655752, -23.8816542884, 57.1497976074, -23.3449664099, -97.5838968887, -60.7349829418};
test_label[706] = '{-4.0143842342};
test_output[706] = '{61.1641818416};
############ END DEBUG ############*/
test_input[5656:5663] = '{32'h41694e24, 32'hc225a1bd, 32'h4091fe09, 32'h3f163993, 32'h41d0f7cd, 32'hc2b77704, 32'hc2981da3, 32'hc2a0cf00};
test_label[707] = '{32'hc2981da3};
test_output[707] = '{32'h42cc5b97};
/*############ DEBUG ############
test_input[5656:5663] = '{14.5815771353, -41.407947142, 4.56226001511, 0.586816030119, 26.1209973879, -91.7324493711, -76.0578820713, -80.404299499};
test_label[707] = '{-76.0578820713};
test_output[707] = '{102.178889198};
############ END DEBUG ############*/
test_input[5664:5671] = '{32'h416c32c4, 32'h4287f7f4, 32'hc26e111d, 32'hc003023a, 32'h4289163a, 32'hc24d2af1, 32'h4275a733, 32'hc1e66527};
test_label[708] = '{32'hc26e111d};
test_output[708] = '{32'h43008347};
/*############ DEBUG ############
test_input[5664:5671] = '{14.7623937101, 67.9842825701, -59.5167121261, -2.04701078493, 68.543413049, -51.291933233, 61.4132820863, -28.7993907036};
test_label[708] = '{-59.5167121261};
test_output[708] = '{128.512796064};
############ END DEBUG ############*/
test_input[5672:5679] = '{32'hc1e7172f, 32'h4299678e, 32'hc2a76e7e, 32'h42b97336, 32'hc1fa58bd, 32'hc2aa9eb8, 32'hc0b1dc03, 32'h4284549c};
test_label[709] = '{32'h4299678e};
test_output[709] = '{32'h41802e9f};
/*############ DEBUG ############
test_input[5672:5679] = '{-28.8863203922, 76.7022588305, -83.7158079186, 92.7250232877, -31.2933293296, -85.3099999187, -5.55810703879, 66.1652512436};
test_label[709] = '{76.7022588305};
test_output[709] = '{16.0227645673};
############ END DEBUG ############*/
test_input[5680:5687] = '{32'h423bcff6, 32'hc297a544, 32'h40c548ad, 32'h423cd721, 32'h4283f167, 32'hc1c3fcca, 32'h42365d8e, 32'hc2783793};
test_label[710] = '{32'hc1c3fcca};
test_output[710] = '{32'h42b4f09a};
/*############ DEBUG ############
test_input[5680:5687] = '{46.9530887383, -75.8227812305, 6.16512139162, 47.210088627, 65.9714908081, -24.4984319606, 45.5913620401, -62.0542724266};
test_label[710] = '{-24.4984319606};
test_output[710] = '{90.4699227827};
############ END DEBUG ############*/
test_input[5688:5695] = '{32'hc213a4c6, 32'h429d618e, 32'hc1c497d3, 32'hc298aeab, 32'hc1bb380b, 32'h4177db42, 32'hc2be2ec5, 32'hc2b8db37};
test_label[711] = '{32'hc213a4c6};
test_output[711] = '{32'h42e733f2};
/*############ DEBUG ############
test_input[5688:5695] = '{-36.9109123568, 78.6905398393, -24.5741319872, -76.3411505972, -23.4023642877, 15.4910294602, -95.0913461997, -92.4281547765};
test_label[711] = '{-36.9109123568};
test_output[711] = '{115.601452196};
############ END DEBUG ############*/
test_input[5696:5703] = '{32'hc106003d, 32'h4293762b, 32'hc261897b, 32'hc2b5e2fb, 32'h40ff9156, 32'h3ecc34a3, 32'hc29e61e5, 32'hc18d0b64};
test_label[712] = '{32'hc2b5e2fb};
test_output[712] = '{32'h4324ac93};
/*############ DEBUG ############
test_input[5696:5703] = '{-8.37505859963, 73.73079827, -56.3842589251, -90.9433242469, 7.98649129265, 0.398839097411, -79.1912040117, -17.6305626958};
test_label[712] = '{-90.9433242469};
test_output[712] = '{164.674122517};
############ END DEBUG ############*/
test_input[5704:5711] = '{32'hc16662f2, 32'hc2902917, 32'h4201c838, 32'h3fa575cf, 32'h4291eb93, 32'hbede5205, 32'h42a4707c, 32'h42376fdf};
test_label[713] = '{32'h4291eb93};
test_output[713] = '{32'h411427a8};
/*############ DEBUG ############
test_input[5704:5711] = '{-14.3991569246, -72.0802573894, 32.4455258044, 1.29265776763, 72.9601091707, -0.434219507976, 82.2196952363, 45.8592489645};
test_label[713] = '{72.9601091707};
test_output[713] = '{9.25968125584};
############ END DEBUG ############*/
test_input[5712:5719] = '{32'h42af34d7, 32'h42404783, 32'hc14a48e2, 32'hc1ea3c43, 32'hc10023d7, 32'hc1fea955, 32'hc2b02516, 32'hc1b2633e};
test_label[714] = '{32'hc1ea3c43};
test_output[714] = '{32'h42e9c3e8};
/*############ DEBUG ############
test_input[5712:5719] = '{87.6032050286, 48.0698361374, -12.6427933077, -29.2794249833, -8.00874980373, -31.8326819584, -88.0724330868, -22.2984585015};
test_label[714] = '{-29.2794249833};
test_output[714] = '{116.882630012};
############ END DEBUG ############*/
test_input[5720:5727] = '{32'h41bb3277, 32'hc28cb6a8, 32'h42c06a71, 32'hc1e2a63f, 32'h42986a69, 32'hc2140882, 32'hc2b92615, 32'h420970e8};
test_label[715] = '{32'hc2b92615};
test_output[715] = '{32'h433cc843};
/*############ DEBUG ############
test_input[5720:5727] = '{23.3996411977, -70.3567526098, 96.2078927792, -28.3311752553, 76.2078328604, -37.0083098888, -92.574378728, 34.3602587194};
test_label[715] = '{-92.574378728};
test_output[715] = '{188.782271509};
############ END DEBUG ############*/
test_input[5728:5735] = '{32'hc2976f84, 32'hc1cf6b0a, 32'hc2a35da1, 32'h4075e4bd, 32'h4199f568, 32'h418c5f57, 32'h416f157b, 32'h4282f8d9};
test_label[716] = '{32'hc2976f84};
test_output[716] = '{32'h430d342e};
/*############ DEBUG ############
test_input[5728:5735] = '{-75.7178037047, -25.9272657542, -81.6828670028, 3.84208599482, 19.2448273314, 17.5465520799, 14.9427441305, 65.4860300343};
test_label[716] = '{-75.7178037047};
test_output[716] = '{141.203833739};
############ END DEBUG ############*/
test_input[5736:5743] = '{32'hc18760a7, 32'hc07edccd, 32'h42848f4d, 32'hc1d82d86, 32'h42bedb96, 32'hc2af86e0, 32'hc2bc1a35, 32'h41be6b67};
test_label[717] = '{32'h42848f4d};
test_output[717] = '{32'h41e93124};
/*############ DEBUG ############
test_input[5736:5743] = '{-16.9221928159, -3.98222657039, 66.2798873822, -27.0222278224, 95.4288822938, -87.7634303429, -94.051182234, 23.802443153};
test_label[717] = '{66.2798873822};
test_output[717] = '{29.1489949116};
############ END DEBUG ############*/
test_input[5744:5751] = '{32'h4230ef24, 32'h4297a34f, 32'hc1c3c314, 32'h42892a2a, 32'hc28d8e55, 32'h428edaa6, 32'hc282eec9, 32'hc200a742};
test_label[718] = '{32'hc1c3c314};
test_output[718] = '{32'h42c89abe};
/*############ DEBUG ############
test_input[5744:5751] = '{44.2335343992, 75.8189619644, -24.4702538791, 68.5823541822, -70.7779902316, 71.4270511536, -65.4663784675, -32.1633363687};
test_label[718] = '{-24.4702538791};
test_output[718] = '{100.302227627};
############ END DEBUG ############*/
test_input[5752:5759] = '{32'hc2aead47, 32'h42a98a97, 32'h424f0a04, 32'h423a199e, 32'hc22bc21e, 32'h3fb96581, 32'h41576262, 32'h40458ce1};
test_label[719] = '{32'h41576262};
test_output[719] = '{32'h428e9e4b};
/*############ DEBUG ############
test_input[5752:5759] = '{-87.3384359554, 84.7706817244, 51.7597815703, 46.5250149708, -42.9395691224, 1.44841016288, 13.4615189793, 3.08672349611};
test_label[719] = '{13.4615189793};
test_output[719] = '{71.3091627451};
############ END DEBUG ############*/
test_input[5760:5767] = '{32'hc288d814, 32'h424f91dd, 32'hc267dca7, 32'hc0c0291c, 32'h42815ddd, 32'h424e382f, 32'hc2c23c22, 32'hc15cf253};
test_label[720] = '{32'hc288d814};
test_output[720] = '{32'h43051af9};
/*############ DEBUG ############
test_input[5760:5767] = '{-68.4220266078, 51.8924457215, -57.9654793679, -6.00501844013, 64.6833282002, 51.5548682604, -97.1174454115, -13.8091607825};
test_label[720] = '{-68.4220266078};
test_output[720] = '{133.105359582};
############ END DEBUG ############*/
test_input[5768:5775] = '{32'h41ce2342, 32'hc0d17568, 32'hc19718c2, 32'h42bb498b, 32'hc2a34424, 32'hc2b1129d, 32'hc10250f0, 32'hc27d6f24};
test_label[721] = '{32'hc10250f0};
test_output[721] = '{32'h42cb93a9};
/*############ DEBUG ############
test_input[5768:5775] = '{25.7672150415, -6.54558187245, -18.8870890769, 93.6436353957, -81.6330892438, -88.5363571628, -8.14475979192, -63.3585360055};
test_label[721] = '{-8.14475979192};
test_output[721] = '{101.788395188};
############ END DEBUG ############*/
test_input[5776:5783] = '{32'h41ec372c, 32'hc1026d75, 32'h428c0083, 32'hc2ac5e61, 32'h4241a149, 32'h429b253d, 32'hc2b72663, 32'hc22c327d};
test_label[722] = '{32'h428c0083};
test_output[722] = '{32'h40f24fd3};
/*############ DEBUG ############
test_input[5776:5783] = '{29.5269403306, -8.15172300635, 70.0009983692, -86.1843346113, 48.4075059911, 77.572727963, -91.5749771273, -43.0493046361};
test_label[722] = '{70.0009983692};
test_output[722] = '{7.57224426267};
############ END DEBUG ############*/
test_input[5784:5791] = '{32'hc28bcfd2, 32'hc1c3bfe0, 32'hc2b1c2b1, 32'hc23e250e, 32'h428a4192, 32'hc2a1f623, 32'hc229561d, 32'hc2599ec2};
test_label[723] = '{32'hc28bcfd2};
test_output[723] = '{32'h430b08b2};
/*############ DEBUG ############
test_input[5784:5791] = '{-69.9059028163, -24.4686897782, -88.8802582643, -47.5361862781, 69.128066153, -80.9807338577, -42.3340968381, -54.4050382802};
test_label[723] = '{-69.9059028163};
test_output[723] = '{139.033968969};
############ END DEBUG ############*/
test_input[5792:5799] = '{32'hc2c2660f, 32'h41909d75, 32'hc29af0fe, 32'hc2a46175, 32'hc2a9f16d, 32'hc2366c0d, 32'hc22815a6, 32'hc29f409e};
test_label[724] = '{32'hc2366c0d};
test_output[724] = '{32'h427ebac7};
/*############ DEBUG ############
test_input[5792:5799] = '{-97.1993339307, 18.0768835474, -77.4706894543, -82.1903464818, -84.9715377084, -45.6055173363, -42.0211418955, -79.6262082973};
test_label[724] = '{-45.6055173363};
test_output[724] = '{63.6824008837};
############ END DEBUG ############*/
test_input[5800:5807] = '{32'h4242d7c8, 32'hc1ed70be, 32'hc14a37cb, 32'h420e6dcb, 32'h4234fece, 32'h42a93fd6, 32'hc1e5d62f, 32'h40439672};
test_label[725] = '{32'h4242d7c8};
test_output[725] = '{32'h420fa7e3};
/*############ DEBUG ############
test_input[5800:5807] = '{48.7107243459, -29.6800496897, -12.6386214371, 35.6072180934, 45.2488308215, 84.624677172, -28.7295816708, 3.05605737843};
test_label[725] = '{48.7107243459};
test_output[725] = '{35.913952826};
############ END DEBUG ############*/
test_input[5808:5815] = '{32'h4268ef20, 32'hc2bee713, 32'h3d96d996, 32'hc1202669, 32'hc0f0fdaa, 32'h428f3e58, 32'hc2579e43, 32'hc1e42a87};
test_label[726] = '{32'hc1e42a87};
test_output[726] = '{32'h42c848fa};
/*############ DEBUG ############
test_input[5808:5815] = '{58.2335191006, -95.4513156254, 0.0736571984036, -10.009377135, -7.53096504372, 71.6217683481, -53.9045519022, -28.5207648751};
test_label[726] = '{-28.5207648751};
test_output[726] = '{100.142534756};
############ END DEBUG ############*/
test_input[5816:5823] = '{32'h4145f383, 32'hc292de52, 32'hc2790f73, 32'h429ad60a, 32'h41ad026a, 32'hc2a14b2d, 32'hc202466a, 32'hc2665ed4};
test_label[727] = '{32'h429ad60a};
test_output[727] = '{32'h80000000};
/*############ DEBUG ############
test_input[5816:5823] = '{12.3719513451, -73.4342203845, -62.2650884239, 77.4180421841, 21.6261792389, -80.6468312658, -32.5687618556, -57.5926045434};
test_label[727] = '{77.4180421841};
test_output[727] = '{-0.0};
############ END DEBUG ############*/
test_input[5824:5831] = '{32'hc1beda28, 32'hc27e6657, 32'h4233b433, 32'h4230ff1b, 32'hc0573c83, 32'h41ca8747, 32'h418c033d, 32'hbf03288c};
test_label[728] = '{32'hc1beda28};
test_output[728] = '{32'h428a6309};
/*############ DEBUG ############
test_input[5824:5831] = '{-23.8565211031, -63.5999425295, 44.9259753152, 44.2491277337, -3.36306836572, 25.3160528421, 17.5015820221, -0.512337428239};
test_label[728] = '{-23.8565211031};
test_output[728] = '{69.1934243011};
############ END DEBUG ############*/
test_input[5832:5839] = '{32'hc2695177, 32'h42584d6b, 32'h42c736b5, 32'hc2143111, 32'hc24e44fb, 32'h40c7b8ea, 32'hc2bc8a59, 32'h42a985d9};
test_label[729] = '{32'hc2143111};
test_output[729] = '{32'h4308a79f};
/*############ DEBUG ############
test_input[5832:5839] = '{-58.3295540216, 54.0756017702, 99.6068479303, -37.0479152404, -51.5673618751, 6.24132261424, -94.2702098091, 84.7614238657};
test_label[729] = '{-37.0479152404};
test_output[729] = '{136.654763528};
############ END DEBUG ############*/
test_input[5840:5847] = '{32'h42ab6a74, 32'h42ace95c, 32'h42077c2b, 32'h42945375, 32'h42374902, 32'hc20af00a, 32'hc18b567a, 32'hc143a03a};
test_label[730] = '{32'h42ace95c};
test_output[730] = '{32'h3ec66e6a};
/*############ DEBUG ############
test_input[5840:5847] = '{85.7079164758, 86.4557765807, 33.8712572744, 74.1629985793, 45.8212969727, -34.734412483, -17.4172241611, -12.2266175334};
test_label[730] = '{86.4557765807};
test_output[730] = '{0.387561140776};
############ END DEBUG ############*/
test_input[5848:5855] = '{32'hc2984a3f, 32'hc1ab7847, 32'h420407c0, 32'hc26265bf, 32'h42800c0b, 32'hc236bccc, 32'hc21c2f35, 32'hc1b92d88};
test_label[731] = '{32'hc236bccc};
test_output[731] = '{32'h42db6a71};
/*############ DEBUG ############
test_input[5848:5855] = '{-76.1450099929, -21.4337283764, 33.0075665962, -56.5993617156, 64.0235237294, -45.6843707588, -39.0461024363, -23.1472316884};
test_label[731] = '{-45.6843707588};
test_output[731] = '{109.707894488};
############ END DEBUG ############*/
test_input[5856:5863] = '{32'h4280b70f, 32'h426494e4, 32'h42b8834d, 32'hc29a5658, 32'h42ad0d72, 32'hc257a05a, 32'hc2973279, 32'h42ac4756};
test_label[732] = '{32'h42ac4756};
test_output[732] = '{32'h40c3ebff};
/*############ DEBUG ############
test_input[5856:5863] = '{64.3575351279, 57.1453992191, 92.2564468451, -77.1686390897, 86.5262614897, -53.9065936715, -75.5985831845, 86.1393250569};
test_label[732] = '{86.1393250569};
test_output[732] = '{6.12255825196};
############ END DEBUG ############*/
test_input[5864:5871] = '{32'h4230ad0b, 32'hc020f709, 32'hc279f2ff, 32'hc1d56508, 32'h42aa6108, 32'h42a33ed2, 32'hc2ad9c8e, 32'h42093bac};
test_label[733] = '{32'hc2ad9c8e};
test_output[733] = '{32'h432c05ed};
/*############ DEBUG ############
test_input[5864:5871] = '{44.1689864924, -2.51507791852, -62.4872999765, -26.6743311903, 85.1895170223, 81.6226970942, -86.8057737783, 34.3082728833};
test_label[733] = '{-86.8057737783};
test_output[733] = '{172.023144785};
############ END DEBUG ############*/
test_input[5872:5879] = '{32'hc2a40e99, 32'h4275d187, 32'hc29baa8b, 32'h424e6583, 32'hbed9a869, 32'hc0b53f10, 32'h41661b41, 32'h40613242};
test_label[734] = '{32'h41661b41};
test_output[734] = '{32'h423c4ac5};
/*############ DEBUG ############
test_input[5872:5879] = '{-82.0285074491, 61.4546170961, -77.8330918299, 51.5991315841, -0.425112977738, -5.66394810139, 14.3816540109, 3.51869256581};
test_label[734] = '{14.3816540109};
test_output[734] = '{47.0730155424};
############ END DEBUG ############*/
test_input[5880:5887] = '{32'hc2901526, 32'hc291ae58, 32'h4221848d, 32'h429a4b7a, 32'hc25da26d, 32'hc286e78d, 32'h4275ea18, 32'h416d2e9a};
test_label[735] = '{32'h429a4b7a};
test_output[735] = '{32'h342846b4};
/*############ DEBUG ############
test_input[5880:5887] = '{-72.0413073658, -72.8405129206, 40.3794458988, 77.147417389, -55.4086197638, -67.4522466867, 61.4786085947, 14.823877461};
test_label[735] = '{77.147417389};
test_output[735] = '{1.5671940319e-07};
############ END DEBUG ############*/
test_input[5888:5895] = '{32'hc08f9e59, 32'h4222b1ed, 32'hc2c79add, 32'h421dc204, 32'hc2375532, 32'hc2225104, 32'h428e88d0, 32'hc2bb0102};
test_label[736] = '{32'hc08f9e59};
test_output[736] = '{32'h429782b5};
/*############ DEBUG ############
test_input[5888:5895] = '{-4.48807940734, 40.6737551378, -99.8024684103, 39.4394689942, -45.83319716, -40.5791180812, 71.2672114038, -93.5019663601};
test_label[736] = '{-4.48807940734};
test_output[736] = '{75.7552908111};
############ END DEBUG ############*/
test_input[5896:5903] = '{32'hc299aae5, 32'h428239d2, 32'hc2669fbe, 32'hc1bb5185, 32'h41a3120b, 32'h4221ee53, 32'hc21c1810, 32'h42c0661a};
test_label[737] = '{32'hc2669fbe};
test_output[737] = '{32'h4319dafc};
/*############ DEBUG ############
test_input[5896:5903] = '{-76.8337813407, 65.112933001, -57.6559965265, -23.4148046298, 20.3838107204, 40.4827394705, -39.0234974512, 96.1994172257};
test_label[737] = '{-57.6559965265};
test_output[737] = '{153.855413752};
############ END DEBUG ############*/
test_input[5904:5911] = '{32'h41d8afa9, 32'hc1fbba48, 32'h4199c875, 32'hc29edb4f, 32'h41d7187e, 32'hc2188a22, 32'h42930599, 32'hc00da405};
test_label[738] = '{32'hc00da405};
test_output[738] = '{32'h429772b9};
/*############ DEBUG ############
test_input[5904:5911] = '{27.08577065, -31.4659579988, 19.2228792342, -79.4283406284, 26.8869590085, -38.1348969071, 73.5109353859, -2.21313592468};
test_label[738] = '{-2.21313592468};
test_output[738] = '{75.7240713106};
############ END DEBUG ############*/
test_input[5912:5919] = '{32'hc2a4d0f5, 32'h40e3c3a6, 32'hc19e89f4, 32'hc296620f, 32'h42290f2d, 32'hc2235a0c, 32'hc2007523, 32'hc2bc4ba0};
test_label[739] = '{32'h40e3c3a6};
test_output[739] = '{32'h420c96b8};
/*############ DEBUG ############
test_input[5912:5919] = '{-82.4081182823, 7.11763303567, -19.8173602238, -75.1915182962, 42.2648201114, -40.8379357426, -32.1143914183, -94.147707162};
test_label[739] = '{7.11763303567};
test_output[739] = '{35.1471870757};
############ END DEBUG ############*/
test_input[5920:5927] = '{32'h42860ccc, 32'h42bacf19, 32'h41f738de, 32'h425db763, 32'hc19e4925, 32'h424e12c5, 32'hc23c3300, 32'hc25b86b4};
test_label[740] = '{32'h42bacf19};
test_output[740] = '{32'h2c75fe00};
/*############ DEBUG ############
test_input[5920:5927] = '{67.0249967282, 93.4044885457, 30.9027669919, 55.4290874246, -19.7857147379, 51.5183286877, -47.0498063424, -54.8815475202};
test_label[740] = '{93.4044885457};
test_output[740] = '{3.49575923764e-12};
############ END DEBUG ############*/
test_input[5928:5935] = '{32'hc22e8509, 32'hc1fc4d66, 32'h427399a2, 32'h41dc8139, 32'hc28efb25, 32'h40f913cb, 32'h41c2cb46, 32'hc15dcfaf};
test_label[741] = '{32'h41dc8139};
test_output[741] = '{32'h42055906};
/*############ DEBUG ############
test_input[5928:5935] = '{-43.6299169441, -31.5377925929, 60.9000334899, 27.5630978792, -71.4905180425, 7.78366617166, 24.3492552836, -13.8632036179};
test_label[741] = '{27.5630978792};
test_output[741] = '{33.3369356107};
############ END DEBUG ############*/
test_input[5936:5943] = '{32'hc2440faa, 32'hc1ca8b93, 32'hc0e68693, 32'hc2b66659, 32'hc1d7b2cf, 32'hbf1ba1f7, 32'hc1e78d2c, 32'hc2b4535f};
test_label[742] = '{32'hc1ca8b93};
test_output[742] = '{32'h41c5b14f};
/*############ DEBUG ############
test_input[5936:5943] = '{-49.0152985507, -25.3181521613, -7.20392747989, -91.1999013418, -26.9623080974, -0.607940149708, -28.9439309878, -90.1628374818};
test_label[742] = '{-25.3181521613};
test_output[742] = '{24.7115769174};
############ END DEBUG ############*/
test_input[5944:5951] = '{32'h42b8bc5f, 32'hc29fefc3, 32'h4211700a, 32'h4150e69d, 32'h42143425, 32'h41905dcd, 32'h40cb334a, 32'hc248e52c};
test_label[743] = '{32'h41905dcd};
test_output[743] = '{32'h4294a4eb};
/*############ DEBUG ############
test_input[5944:5951] = '{92.367910709, -79.9682868077, 36.3594136282, 13.0563016922, 37.0509230567, 18.0458017119, 6.35001076407, -50.2237998453};
test_label[743] = '{18.0458017119};
test_output[743] = '{74.3221089971};
############ END DEBUG ############*/
test_input[5952:5959] = '{32'hc28d550d, 32'hc2a58d67, 32'h424084a6, 32'h3e2e3c16, 32'hc2adc319, 32'h41e3e8bd, 32'hc2bb4887, 32'h417971cd};
test_label[744] = '{32'h41e3e8bd};
test_output[744] = '{32'h419d208e};
/*############ DEBUG ############
test_input[5952:5959] = '{-70.6661137959, -82.7761742936, 48.1295377442, 0.170151077729, -86.88104949, 28.4886416069, -93.6416557594, 15.5902834005};
test_label[744] = '{28.4886416069};
test_output[744] = '{19.6408961402};
############ END DEBUG ############*/
test_input[5960:5967] = '{32'h4260176f, 32'hc2c20cc0, 32'h4203ba35, 32'h42552ac0, 32'hc2bd4331, 32'h4206df74, 32'hc2aa38a0, 32'hc22b6249};
test_label[745] = '{32'hc2c20cc0};
test_output[745] = '{32'h43191c64};
/*############ DEBUG ############
test_input[5960:5967] = '{56.0228855662, -97.0249059371, 32.9318441198, 53.2917494829, -94.6312324524, 33.7182175189, -85.1105961326, -42.8459801201};
test_label[745] = '{-97.0249059371};
test_output[745] = '{153.110902666};
############ END DEBUG ############*/
test_input[5968:5975] = '{32'hc249d7c5, 32'h428a612d, 32'h42a19f76, 32'hc1b69e1a, 32'hc2794bc1, 32'hc22ab7e7, 32'hc2a17541, 32'hc234ff85};
test_label[746] = '{32'h42a19f76};
test_output[746] = '{32'h37167c9f};
/*############ DEBUG ############
test_input[5968:5975] = '{-50.4607130614, 69.1897949838, 80.8114474465, -22.8271972819, -62.3239779677, -42.6795934255, -80.7290094696, -45.2495291053};
test_label[746] = '{80.8114474465};
test_output[746] = '{8.96971237545e-06};
############ END DEBUG ############*/
test_input[5976:5983] = '{32'h41599766, 32'hc02cdd4f, 32'h42386a9f, 32'h42b2e419, 32'h419ea15b, 32'hc026a0b5, 32'h42ada3c1, 32'hc1786905};
test_label[747] = '{32'h42b2e419};
test_output[747] = '{32'h3d8f22ea};
/*############ DEBUG ############
test_input[5976:5983] = '{13.5994623761, -2.70100758486, 46.104121946, 89.4455058723, 19.828787411, -2.60355887795, 86.8198336976, -15.5256398189};
test_label[747] = '{89.4455058723};
test_output[747] = '{0.0698908106961};
############ END DEBUG ############*/
test_input[5984:5991] = '{32'hc2836706, 32'hc20afb65, 32'h428f30a7, 32'hc155cb31, 32'hc175cba4, 32'h42a10fbb, 32'h41d2d694, 32'h40e0b3b5};
test_label[748] = '{32'h428f30a7};
test_output[748] = '{32'h410ef928};
/*############ DEBUG ############
test_input[5984:5991] = '{-65.7012167277, -34.7455036583, 71.5950237579, -13.362107571, -15.3622167818, 80.5307213318, 26.3547735695, 7.02193705528};
test_label[748] = '{71.5950237579};
test_output[748] = '{8.93582917126};
############ END DEBUG ############*/
test_input[5992:5999] = '{32'h422e38cb, 32'hc29ef34a, 32'hc1e7a6b8, 32'h42904ddd, 32'hc16044f2, 32'h428fbd57, 32'hc1401d2e, 32'hc1621783};
test_label[749] = '{32'h428fbd57};
test_output[749] = '{32'h3f581e20};
/*############ DEBUG ############
test_input[5992:5999] = '{43.5554622308, -79.4751732766, -28.9564061043, 72.1520739484, -14.0168324751, 71.8698024724, -12.0071242074, -14.1307399834};
test_label[749] = '{71.8698024724};
test_output[749] = '{0.844209676495};
############ END DEBUG ############*/
test_input[6000:6007] = '{32'hc20b1d76, 32'hc20f4eb7, 32'hc21a2d1a, 32'hc2a1d01d, 32'hc2295d8d, 32'hc2452588, 32'hc2574c8f, 32'h4209464e};
test_label[750] = '{32'hc2295d8d};
test_output[750] = '{32'h429951ed};
/*############ DEBUG ############
test_input[6000:6007] = '{-34.7787692338, -35.826869562, -38.5440448446, -80.9064718997, -42.3413570722, -49.2866523899, -53.824764638, 34.3186575329};
test_label[750] = '{-42.3413570722};
test_output[750] = '{76.6600146051};
############ END DEBUG ############*/
test_input[6008:6015] = '{32'h41d172e1, 32'h419c040c, 32'hc2b7a329, 32'h411a0e12, 32'h41904f11, 32'h40280c04, 32'h3ff17016, 32'h42b89d81};
test_label[751] = '{32'h3ff17016};
test_output[751] = '{32'h42b4d7c1};
/*############ DEBUG ############
test_input[6008:6015] = '{26.1810930849, 19.5019765333, -91.8186725663, 9.62843525101, 18.0386066312, 2.6257334075, 1.8862330825, 92.3076250965};
test_label[751] = '{1.8862330825};
test_output[751] = '{90.421392014};
############ END DEBUG ############*/
test_input[6016:6023] = '{32'h428892c7, 32'h42b4f29b, 32'h42617e0e, 32'hc28b5385, 32'hc2303d6c, 32'hc1fed953, 32'h4218fad2, 32'h4215b937};
test_label[752] = '{32'h4218fad2};
test_output[752] = '{32'h4250ea65};
/*############ DEBUG ############
test_input[6016:6023] = '{68.2866766178, 90.4738407576, 56.3731006613, -69.6631231373, -44.0599834851, -31.8561147529, 38.244941203, 37.4308757142};
test_label[752] = '{38.244941203};
test_output[752] = '{52.2288995548};
############ END DEBUG ############*/
test_input[6024:6031] = '{32'h42abf9d0, 32'h428794cf, 32'hc24c1357, 32'hc19210a8, 32'h421f7c92, 32'h42b63c1e, 32'h42659421, 32'h3f734f94};
test_label[753] = '{32'h42659421};
test_output[753] = '{32'h4206ea27};
/*############ DEBUG ############
test_input[6024:6031] = '{85.9879116701, 67.7906390604, -51.0188848189, -18.2581335295, 39.8716520044, 91.1174200213, 57.3946581079, 0.950433010348};
test_label[753] = '{57.3946581079};
test_output[753] = '{33.7286639323};
############ END DEBUG ############*/
test_input[6032:6039] = '{32'h42539a8c, 32'h42bf14f1, 32'hc295ae54, 32'hc235d6c4, 32'h424179cb, 32'hc1a6b207, 32'hc2a7f6a8, 32'h424abb13};
test_label[754] = '{32'hc295ae54};
test_output[754] = '{32'h432a61a3};
/*############ DEBUG ############
test_input[6032:6039] = '{52.9009264824, 95.5409007105, -74.8404874349, -45.4597312928, 48.368936677, -20.8369265124, -83.9817467553, 50.6826877607};
test_label[754] = '{-74.8404874349};
test_output[754] = '{170.381388145};
############ END DEBUG ############*/
test_input[6040:6047] = '{32'hc1af4e21, 32'hc151b5da, 32'h42c15138, 32'hc20844a3, 32'h428eab7b, 32'h3fb9d8ef, 32'hc1895ed3, 32'hc2af8149};
test_label[755] = '{32'hc151b5da};
test_output[755] = '{32'h42db87f4};
/*############ DEBUG ############
test_input[6040:6047] = '{-21.913149409, -13.106897004, 96.6586338826, -34.0670289442, 71.3349251082, 1.4519327719, -17.1713004695, -87.7525125798};
test_label[755] = '{-13.106897004};
test_output[755] = '{109.765530887};
############ END DEBUG ############*/
test_input[6048:6055] = '{32'h3fab8b36, 32'hc2a1a40c, 32'hc2bbdbea, 32'h42c6b8c8, 32'hc19c8fd7, 32'h428dab3d, 32'h42b798cc, 32'h42b96dc9};
test_label[756] = '{32'h42b96dc9};
test_output[756] = '{32'h40d4bed9};
/*############ DEBUG ############
test_input[6048:6055] = '{1.34018587842, -80.8204018091, -93.9295191129, 99.360902161, -19.5702336317, 70.8344480289, 91.7984307817, 92.7144217935};
test_label[756] = '{92.7144217935};
test_output[756] = '{6.64829689085};
############ END DEBUG ############*/
test_input[6056:6063] = '{32'h419357e1, 32'hc2689d04, 32'h428a056b, 32'hc24e38b4, 32'h40eabcb8, 32'h4209c38e, 32'h42623436, 32'h42950006};
test_label[757] = '{32'h428a056b};
test_output[757] = '{32'h40afcb69};
/*############ DEBUG ############
test_input[6056:6063] = '{18.4179090063, -58.1533369124, 69.0105833111, -51.5553751676, 7.33553693959, 34.4409730334, 56.5509861278, 74.5000422197};
test_label[757] = '{69.0105833111};
test_output[757] = '{5.4935804976};
############ END DEBUG ############*/
test_input[6064:6071] = '{32'h409e071c, 32'h408780fd, 32'hc2319cda, 32'h429c7919, 32'hc2a01808, 32'h428fc95a, 32'hc22090a3, 32'hc2636a11};
test_label[758] = '{32'h408780fd};
test_output[758] = '{32'h429401ef};
/*############ DEBUG ############
test_input[6064:6071] = '{4.93836786478, 4.23449553084, -44.4031735618, 78.2365182061, -80.0469334352, 71.8932676121, -40.1412450997, -56.8535798196};
test_label[758] = '{4.23449553084};
test_output[758] = '{74.0037797073};
############ END DEBUG ############*/
test_input[6072:6079] = '{32'h409a21f0, 32'hc2a8d24c, 32'h421c8801, 32'h42765f15, 32'h401e3eb7, 32'hc28ddf70, 32'h42b6686b, 32'hc2a6d00a};
test_label[759] = '{32'hc2a8d24c};
test_output[759] = '{32'h432f9d5b};
/*############ DEBUG ############
test_input[6072:6079] = '{4.81664256221, -84.41073612, 39.1328161488, 61.5928554448, 2.4725777153, -70.9364018807, 91.2039403217, -83.4063296419};
test_label[759] = '{-84.41073612};
test_output[759] = '{175.614676442};
############ END DEBUG ############*/
test_input[6080:6087] = '{32'h42896d52, 32'hc272c63e, 32'hc2142b60, 32'hc2a014af, 32'h41019a3f, 32'hc17a03be, 32'hc2845300, 32'h42abb012};
test_label[760] = '{32'h41019a3f};
test_output[760] = '{32'h429b7cca};
/*############ DEBUG ############
test_input[6080:6087] = '{68.7135199596, -60.6935945959, -37.0423586775, -80.040398037, 8.10015759381, -15.6259133553, -66.1621080914, 85.8438870766};
test_label[760] = '{8.10015759381};
test_output[760] = '{77.7437295191};
############ END DEBUG ############*/
test_input[6088:6095] = '{32'hc218c716, 32'h4281a0e2, 32'hc282326b, 32'h4235ff0e, 32'hc2586283, 32'hc2a67706, 32'h41945590, 32'h4294e536};
test_label[761] = '{32'hc2a67706};
test_output[761] = '{32'h431dae22};
/*############ DEBUG ############
test_input[6088:6095] = '{-38.1944210978, 64.8142270851, -65.0984744482, 45.4990758304, -54.0962019316, -83.2324693238, 18.5417784309, 74.4476739659};
test_label[761] = '{-83.2324693238};
test_output[761] = '{157.680208788};
############ END DEBUG ############*/
test_input[6096:6103] = '{32'hc1b3ce88, 32'hc2c72ba7, 32'hc29260cb, 32'h41b57c53, 32'hc20db8a9, 32'hc208697c, 32'h42b2fab6, 32'h428954bd};
test_label[762] = '{32'hc20db8a9};
test_output[762] = '{32'h42f9d70a};
/*############ DEBUG ############
test_input[6096:6103] = '{-22.4758451584, -99.5852577351, -73.1890517934, 22.6857060514, -35.4303323849, -34.103011923, 89.4896682166, 68.6655030637};
test_label[762] = '{-35.4303323849};
test_output[762] = '{124.920000602};
############ END DEBUG ############*/
test_input[6104:6111] = '{32'hc23759e3, 32'hc0d2295f, 32'h401eb2c4, 32'hc29ac470, 32'h3fb8f8ee, 32'h41a309ef, 32'hc1ee9e96, 32'h41fab004};
test_label[763] = '{32'h41a309ef};
test_output[763] = '{32'h412f4c3d};
/*############ DEBUG ############
test_input[6104:6111] = '{-45.8377800635, -6.56755004713, 2.47966087109, -77.3836662164, 1.44509670662, 20.3798497741, -29.8274346962, 31.3359451694};
test_label[763] = '{20.3798497741};
test_output[763] = '{10.9561128464};
############ END DEBUG ############*/
test_input[6112:6119] = '{32'hc2664f76, 32'hc2b09d8d, 32'hc223365b, 32'hc25f7ded, 32'h4297759a, 32'hc2a56214, 32'h4217eb8c, 32'hc2211ab1};
test_label[764] = '{32'hc2664f76};
test_output[764] = '{32'h43054eaa};
/*############ DEBUG ############
test_input[6112:6119] = '{-57.5775981599, -88.307713575, -40.8030818364, -55.8729748146, 75.7296873088, -82.691561407, 37.9800261844, -40.2760670116};
test_label[764] = '{-57.5775981599};
test_output[764] = '{133.307285469};
############ END DEBUG ############*/
test_input[6120:6127] = '{32'h42ba21e2, 32'hc2b3f3d3, 32'h418fb8a2, 32'hc0f94251, 32'h42a10db6, 32'hc24e0173, 32'hc2227631, 32'hc15eb51e};
test_label[765] = '{32'hc24e0173};
test_output[765] = '{32'h4310914e};
/*############ DEBUG ############
test_input[6120:6127] = '{93.0661773578, -89.97621623, 17.9651522735, -7.78934520144, 80.5267758209, -51.5014169674, -40.6154226886, -13.9192183325};
test_label[765] = '{-51.5014169674};
test_output[765] = '{144.567597908};
############ END DEBUG ############*/
test_input[6128:6135] = '{32'h4286bf77, 32'h421007bd, 32'h42a78bbb, 32'h42b1e9de, 32'hc168083a, 32'hc2032638, 32'hc11561d4, 32'h41d950e3};
test_label[766] = '{32'h4286bf77};
test_output[766] = '{32'h41acb50f};
/*############ DEBUG ############
test_input[6128:6135] = '{67.3739514612, 36.0075574557, 83.772913702, 88.9567687168, -14.5020087995, -32.7873231637, -9.33638384197, 27.1644951942};
test_label[766] = '{67.3739514612};
test_output[766] = '{21.5884079511};
############ END DEBUG ############*/
test_input[6136:6143] = '{32'h420f0b58, 32'hc1d351d4, 32'hc2318ffc, 32'hc28bd2e2, 32'h426eac06, 32'hc2be6951, 32'hc23144c4, 32'hc29e8811};
test_label[767] = '{32'hc1d351d4};
test_output[767] = '{32'h42ac2a78};
/*############ DEBUG ############
test_input[6136:6143] = '{35.7610789578, -26.4149560563, -44.3906098764, -69.9118842427, 59.6679928854, -95.2056970977, -44.3171534689, -79.2657566459};
test_label[767] = '{-26.4149560563};
test_output[767] = '{86.0829489418};
############ END DEBUG ############*/
test_input[6144:6151] = '{32'hc2955cb3, 32'hc275609d, 32'h4293fb91, 32'h42aca20b, 32'hc268472d, 32'hc23040ec, 32'hc28f2446, 32'hc23ceeb9};
test_label[768] = '{32'hc268472d};
test_output[768] = '{32'h431062d1};
/*############ DEBUG ############
test_input[6144:6151] = '{-74.6810496787, -61.3443478684, 73.9913423368, 86.3164889805, -58.0695086088, -44.063400741, -71.5708496708, -47.23312716};
test_label[768] = '{-58.0695086088};
test_output[768] = '{144.386002028};
############ END DEBUG ############*/
test_input[6152:6159] = '{32'hc24b9019, 32'h42656693, 32'hc2b109c7, 32'hc092444a, 32'h42bf7504, 32'h41a5f9c1, 32'hc28a70fb, 32'hc24f1ba1};
test_label[769] = '{32'h42bf7504};
test_output[769] = '{32'h80000000};
/*############ DEBUG ############
test_input[6152:6159] = '{-50.8907195234, 57.3501693406, -88.5190979395, -4.57083599662, 95.7285451585, 20.7469502488, -69.2206633544, -51.776980998};
test_label[769] = '{95.7285451585};
test_output[769] = '{-0.0};
############ END DEBUG ############*/
test_input[6160:6167] = '{32'hc088a933, 32'hc2b20749, 32'hc2904075, 32'hc2a7da36, 32'h4255d316, 32'h40626eac, 32'hc07fc974, 32'h426e4c5a};
test_label[770] = '{32'h4255d316};
test_output[770] = '{32'h40c3dc29};
/*############ DEBUG ############
test_input[6160:6167] = '{-4.27065409069, -89.0142256086, -72.1258940723, -83.9261904753, 53.4561379515, 3.53800491972, -3.99667065429, 59.5745635391};
test_label[770] = '{53.4561379515};
test_output[770] = '{6.12062508692};
############ END DEBUG ############*/
test_input[6168:6175] = '{32'h429ec63d, 32'hc1e828de, 32'h41c31f37, 32'h4281d47b, 32'h424c55a7, 32'hc2680909, 32'h3fd8e200, 32'h40dfc208};
test_label[771] = '{32'h3fd8e200};
test_output[771] = '{32'h429b62b5};
/*############ DEBUG ############
test_input[6168:6175] = '{79.3871869538, -29.0199541408, 24.3902425244, 64.9149994229, 51.0836431434, -58.0088244306, 1.69439701248, 6.99243522162};
test_label[771] = '{1.69439701248};
test_output[771] = '{77.6927904599};
############ END DEBUG ############*/
test_input[6176:6183] = '{32'hc24faeb8, 32'hc2b29afd, 32'h42674c08, 32'h41ef7941, 32'hc281829c, 32'h4292b2c1, 32'hc2beed5f, 32'hc2668570};
test_label[772] = '{32'hc2668570};
test_output[772] = '{32'h4302fabc};
/*############ DEBUG ############
test_input[6176:6183] = '{-51.9206248894, -89.3027135315, 57.8242484068, 29.9342061886, -64.7550973301, 73.3491254841, -95.463617818, -57.6303084193};
test_label[772] = '{-57.6303084193};
test_output[772] = '{130.979434084};
############ END DEBUG ############*/
test_input[6184:6191] = '{32'h42a2dc22, 32'h41a9a4ae, 32'hc0fba928, 32'h4199b367, 32'h41e114ae, 32'h42792379, 32'h4180d242, 32'h4211e53e};
test_label[773] = '{32'h41a9a4ae};
test_output[773] = '{32'h4270e5ec};
/*############ DEBUG ############
test_input[6184:6191] = '{81.4299442498, 21.2054096995, -7.86439906833, 19.2125984327, 28.1350983049, 62.2846414584, 16.1026651716, 36.4738705696};
test_label[773] = '{21.2054096995};
test_output[773] = '{60.2245345551};
############ END DEBUG ############*/
test_input[6192:6199] = '{32'hc123e7cd, 32'h41e8f019, 32'h41e50a0e, 32'h42b76aec, 32'h422ece97, 32'h421173b0, 32'hc2393960, 32'hc23c2bba};
test_label[774] = '{32'h41e8f019};
test_output[774] = '{32'h427a5dcc};
/*############ DEBUG ############
test_input[6192:6199] = '{-10.2440922901, 29.1172345922, 28.6299093055, 91.7088338829, 43.7017479242, 36.3629764335, -46.3060307317, -47.0427033146};
test_label[774] = '{29.1172345922};
test_output[774] = '{62.5915992907};
############ END DEBUG ############*/
test_input[6200:6207] = '{32'hc2b398a3, 32'hc1dcbe87, 32'h428f6712, 32'hc12dab0d, 32'h42aab42e, 32'h429bb62a, 32'h42a3f0c4, 32'h42c3b2bb};
test_label[775] = '{32'h42c3b2bb};
test_output[775] = '{32'h3681bb65};
/*############ DEBUG ############
test_input[6200:6207] = '{-89.798118197, -27.593031486, 71.7013090714, -10.8542604061, 85.3519113873, 77.8557918795, 81.9702457249, 97.8490819178};
test_label[775] = '{97.8490819178};
test_output[775] = '{3.86631532695e-06};
############ END DEBUG ############*/
test_input[6208:6215] = '{32'h42bd9afb, 32'h41116391, 32'h4180f0f7, 32'hc2aaa260, 32'h4288bfbb, 32'h42ae3842, 32'h4296cb35, 32'h423dbabf};
test_label[776] = '{32'h4296cb35};
test_output[776] = '{32'h419b4008};
/*############ DEBUG ############
test_input[6208:6215] = '{94.8026951068, 9.08680800625, 16.1176583694, -85.317141876, 68.3744773714, 87.1098800671, 75.3968864296, 47.4323684966};
test_label[776] = '{75.3968864296};
test_output[776] = '{19.4062646694};
############ END DEBUG ############*/
test_input[6216:6223] = '{32'hc24126b4, 32'hc2859447, 32'h42b42bfa, 32'h428372ca, 32'hc2857182, 32'hc262bc3f, 32'hc158a912, 32'h42863c0b};
test_label[777] = '{32'h428372ca};
test_output[777] = '{32'h41c2e4bf};
/*############ DEBUG ############
test_input[6216:6223] = '{-48.2877973896, -66.7896067804, 90.0858908891, 65.7241977864, -66.7216965996, -56.6838347621, -13.541276842, 67.1172688193};
test_label[777] = '{65.7241977864};
test_output[777] = '{24.3616931028};
############ END DEBUG ############*/
test_input[6224:6231] = '{32'hc2685b33, 32'hc26a88bc, 32'h42c1faec, 32'h42a5f086, 32'hc10831a2, 32'hc2024965, 32'hc2b5a555, 32'h42899c87};
test_label[778] = '{32'hc2685b33};
test_output[778] = '{32'h431b1443};
/*############ DEBUG ############
test_input[6224:6231] = '{-58.0890604486, -58.633529848, 96.9900830124, 82.9697687863, -8.51211699756, -32.5716748432, -90.8229166685, 68.8057167836};
test_label[778] = '{-58.0890604486};
test_output[778] = '{155.079144276};
############ END DEBUG ############*/
test_input[6232:6239] = '{32'hc172afd8, 32'h40a26b2f, 32'h4191a9a6, 32'hc2ac8c7c, 32'h42bb1c87, 32'h4203f9e7, 32'h42a29b75, 32'hc2607d0e};
test_label[779] = '{32'h42bb1c87};
test_output[779] = '{32'h36a039f0};
/*############ DEBUG ############
test_input[6232:6239] = '{-15.1679304765, 5.07558410908, 18.20783594, -86.2743848874, 93.5557203066, 32.9940464523, 81.3036304579, -56.1221237705};
test_label[779] = '{93.5557203066};
test_output[779] = '{4.77511626226e-06};
############ END DEBUG ############*/
test_input[6240:6247] = '{32'hc221e6ef, 32'h42abca00, 32'h41e783a9, 32'h425312bb, 32'hc24d0ca2, 32'hc2c2b1db, 32'hc2b82bbf, 32'hc1fd7645};
test_label[780] = '{32'hc2b82bbf};
test_output[780] = '{32'h4331fae0};
/*############ DEBUG ############
test_input[6240:6247] = '{-40.4755217819, 85.8945310001, 28.9392865813, 52.7682919889, -51.2623382616, -97.3473759108, -92.0854428109, -31.6827479548};
test_label[780] = '{-92.0854428109};
test_output[780] = '{177.979973811};
############ END DEBUG ############*/
test_input[6248:6255] = '{32'hc23461ce, 32'h429d69bd, 32'hc025a90b, 32'h4272090d, 32'hc2c0b3b2, 32'hc25b13b9, 32'hc214dc87, 32'hc1e214dc};
test_label[781] = '{32'hc25b13b9};
test_output[781] = '{32'h430579cd};
/*############ DEBUG ############
test_input[6248:6255] = '{-45.0955121769, 78.7065179019, -2.5884424992, 60.5088376747, -96.3509700193, -54.7692609315, -37.215359897, -28.2601860466};
test_label[781] = '{-54.7692609315};
test_output[781] = '{133.475778846};
############ END DEBUG ############*/
test_input[6256:6263] = '{32'hc151e69d, 32'hc2958c8f, 32'hc1c72ba1, 32'hc0c3e911, 32'h424826a7, 32'hc233f76f, 32'hc2a90672, 32'h42c3d90c};
test_label[782] = '{32'hc233f76f};
test_output[782] = '{32'h430eea62};
/*############ DEBUG ############
test_input[6256:6263] = '{-13.1188016181, -74.7745280336, -24.8963026869, -6.12220026144, 50.0377447655, -44.9916328272, -84.5125852671, 97.9239178779};
test_label[782] = '{-44.9916328272};
test_output[782] = '{142.915550705};
############ END DEBUG ############*/
test_input[6264:6271] = '{32'hc140158d, 32'h42351f1c, 32'h416ec0a0, 32'hbff13f93, 32'h41ccdc05, 32'hc2b2e60c, 32'h41dba1e1, 32'h407e60de};
test_label[783] = '{32'h416ec0a0};
test_output[783] = '{32'h41f2dde7};
/*############ DEBUG ############
test_input[6264:6271] = '{-12.0052613173, 45.2803788198, 14.922027672, -1.88475258085, 25.6074323598, -89.4493108147, 27.4540433473, 3.9746623284};
test_label[783] = '{14.922027672};
test_output[783] = '{30.3583511688};
############ END DEBUG ############*/
test_input[6272:6279] = '{32'h3faccce2, 32'hc298a488, 32'hc1521531, 32'hc18c5cb8, 32'h42002136, 32'hc2890ed3, 32'hc27121d2, 32'hc26b3a77};
test_label[784] = '{32'hc1521531};
test_output[784] = '{32'h4234a682};
/*############ DEBUG ############
test_input[6272:6279] = '{1.35000251149, -76.3213487283, -13.1301740425, -17.5452733077, 32.0324312447, -68.5289539236, -60.2830281319, -58.8070929794};
test_label[784] = '{-13.1301740425};
test_output[784] = '{45.1626052872};
############ END DEBUG ############*/
test_input[6280:6287] = '{32'h42006fdf, 32'h42aa211c, 32'h417ac343, 32'hc1c30989, 32'hc2a97ce1, 32'h415d6214, 32'h42527f38, 32'h3d87017e};
test_label[785] = '{32'h417ac343};
test_output[785] = '{32'h428ac8b3};
/*############ DEBUG ############
test_input[6280:6287] = '{32.1092504634, 85.0646651336, 15.6726712198, -24.3796557674, -84.743904351, 13.8364446005, 52.6242366208, 0.0659208115617};
test_label[785] = '{15.6726712198};
test_output[785] = '{69.3919939138};
############ END DEBUG ############*/
test_input[6288:6295] = '{32'h42b01648, 32'hc2b04d86, 32'hc22c594d, 32'h42500d90, 32'h4211896a, 32'hc1a3cba5, 32'hc286d94e, 32'h408be6d8};
test_label[786] = '{32'h408be6d8};
test_output[786] = '{32'h42a757da};
/*############ DEBUG ############
test_input[6288:6295] = '{88.04351426, -88.1514097531, -43.0872066335, 52.0132434846, 36.3841939849, -20.4744351832, -67.4244257375, 4.3719292449};
test_label[786] = '{4.3719292449};
test_output[786] = '{83.6715850151};
############ END DEBUG ############*/
test_input[6296:6303] = '{32'h420fe215, 32'h41acabdf, 32'hc2afb857, 32'hc2aa6743, 32'h425d2022, 32'hc255ca27, 32'hc2b80d2f, 32'h428df6bc};
test_label[787] = '{32'hc255ca27};
test_output[787] = '{32'h42f8dbd0};
/*############ DEBUG ############
test_input[6296:6303] = '{35.9707846512, 21.583921664, -87.8600372497, -85.201686163, 55.2813795278, -53.4474154602, -92.0257491638, 70.9819042451};
test_label[787] = '{-53.4474154602};
test_output[787] = '{124.429319857};
############ END DEBUG ############*/
test_input[6304:6311] = '{32'h42ac94e9, 32'h42a28d53, 32'hc1b87fcf, 32'hc14fce04, 32'hc17b34bb, 32'h422779ad, 32'hc2bac336, 32'h426b3a15};
test_label[788] = '{32'h42a28d53};
test_output[788] = '{32'h40a0af8f};
/*############ DEBUG ############
test_input[6304:6311] = '{86.2908388894, 81.2760254246, -23.0624056255, -12.987797224, -15.700373797, 41.8688227312, -93.3812741296, 58.806720281};
test_label[788] = '{81.2760254246};
test_output[788] = '{5.02143039483};
############ END DEBUG ############*/
test_input[6312:6319] = '{32'h418cfa3b, 32'hc2a2b76e, 32'hc280c8e6, 32'h42c6c0eb, 32'h42c341c6, 32'hc1aa3070, 32'h42264330, 32'h425dcf19};
test_label[789] = '{32'h42c6c0eb};
test_output[789] = '{32'h3e2452b5};
/*############ DEBUG ############
test_input[6312:6319] = '{17.6221835326, -81.3582639898, -64.3923775788, 99.3767935268, 97.6284647676, -21.2736513634, 41.5656110722, 55.4522448402};
test_label[789] = '{99.3767935268};
test_output[789] = '{0.160471749175};
############ END DEBUG ############*/
test_input[6320:6327] = '{32'h427fedec, 32'hc18b2ab7, 32'h4129d5cc, 32'hc1fa4942, 32'hc2b1a5e6, 32'h40a16853, 32'h4297249b, 32'h426a4714};
test_label[790] = '{32'h427fedec};
test_output[790] = '{32'h41396d2f};
/*############ DEBUG ############
test_input[6320:6327] = '{63.9823466062, -17.3958562171, 10.6146960861, -31.2857710172, -88.8240193947, 5.04398474102, 75.5714931594, 58.5694134142};
test_label[790] = '{63.9823466062};
test_output[790] = '{11.5891558606};
############ END DEBUG ############*/
test_input[6328:6335] = '{32'hc0d04e1c, 32'h42a3a797, 32'hc1cada1e, 32'hc2bc429a, 32'hc0b7982b, 32'h420a5fbb, 32'hc2c35142, 32'h42b92e14};
test_label[791] = '{32'h42b92e14};
test_output[791] = '{32'h37b1a11a};
/*############ DEBUG ############
test_input[6328:6335] = '{-6.50953464462, 81.827320541, -25.3565023819, -94.1300803186, -5.73732524218, 34.5934860526, -97.6587098659, 92.589996271};
test_label[791] = '{92.589996271};
test_output[791] = '{2.11750635231e-05};
############ END DEBUG ############*/
test_input[6336:6343] = '{32'hc262db02, 32'hc16614c4, 32'hbd7f6b47, 32'hc24d5a05, 32'h41bb38ba, 32'h428ed9a7, 32'hc1f5f4fa, 32'h429c041b};
test_label[792] = '{32'h41bb38ba};
test_output[792] = '{32'h425a6d44};
/*############ DEBUG ############
test_input[6336:6343] = '{-56.7138743943, -14.380069293, -0.0623581667186, -51.3379116044, 23.4026976247, 71.4251033106, -30.7446180814, 78.0080189521};
test_label[792] = '{23.4026976247};
test_output[792] = '{54.6067041795};
############ END DEBUG ############*/
test_input[6344:6351] = '{32'h4298981e, 32'h4288f947, 32'h42bd33ac, 32'hc2599049, 32'h4143afca, 32'hc2002e48, 32'h426ce3c5, 32'h425e7426};
test_label[793] = '{32'hc2002e48};
test_output[793] = '{32'h42fd4ad0};
/*############ DEBUG ############
test_input[6344:6351] = '{76.2971042694, 68.4868725557, 94.6009243788, -54.3909034207, 12.2304176762, -32.0451971986, 59.2224299991, 55.6134274075};
test_label[793] = '{-32.0451971986};
test_output[793] = '{126.646121589};
############ END DEBUG ############*/
test_input[6352:6359] = '{32'hc2027cb3, 32'hc1e9e834, 32'hbfbf3d3d, 32'h42a1fa36, 32'hc2261cdb, 32'hc28fffa5, 32'h4282cef8, 32'h42c2748e};
test_label[794] = '{32'h42a1fa36};
test_output[794] = '{32'h4181e961};
/*############ DEBUG ############
test_input[6352:6359] = '{-32.6217755133, -29.2383803828, -1.49405638127, 80.988692267, -41.5281783757, -71.9993039259, 65.4042321815, 97.2276476273};
test_label[794] = '{80.988692267};
test_output[794] = '{16.2389554489};
############ END DEBUG ############*/
test_input[6360:6367] = '{32'hc2a35a21, 32'hc1c0d639, 32'hc238a5c2, 32'hc19ebc77, 32'h42778442, 32'h4276f309, 32'h42020015, 32'h4202f60c};
test_label[795] = '{32'h4202f60c};
test_output[795] = '{32'h41ee1be9};
/*############ DEBUG ############
test_input[6360:6367] = '{-81.6760300846, -24.1046011073, -46.161871454, -19.8420238862, 61.8791588039, 61.7373385547, 32.50008166, 32.7402793037};
test_label[795] = '{32.7402793037};
test_output[795] = '{29.7636285749};
############ END DEBUG ############*/
test_input[6368:6375] = '{32'hc136199c, 32'h4183763a, 32'hc1229b7e, 32'h42b29882, 32'h423eaf47, 32'h428c6c95, 32'h426a92f3, 32'hc26915c3};
test_label[796] = '{32'hc1229b7e};
test_output[796] = '{32'h42c6ebf2};
/*############ DEBUG ############
test_input[6368:6375] = '{-11.3812523254, 16.4327274673, -10.1629618438, 89.2978701267, 47.6711701036, 70.2120750448, 58.643504225, -58.2712507918};
test_label[796] = '{-10.1629618438};
test_output[796] = '{99.4608319756};
############ END DEBUG ############*/
test_input[6376:6383] = '{32'h41be16dc, 32'hc2b9e67b, 32'hc29d13da, 32'hc1f25ef0, 32'hc2156c50, 32'h42925482, 32'hc2255045, 32'h41d3f324};
test_label[797] = '{32'hc1f25ef0};
test_output[797] = '{32'h42ceec3e};
/*############ DEBUG ############
test_input[6376:6383] = '{23.7611624585, -92.950158069, -78.5387732453, -30.2963563214, -37.3557744773, 73.1650522461, -41.3283896029, 26.4937209939};
test_label[797] = '{-30.2963563214};
test_output[797] = '{103.461408567};
############ END DEBUG ############*/
test_input[6384:6391] = '{32'h41922e3b, 32'h41ef7585, 32'h418b4ee3, 32'h428ad580, 32'hc2049c76, 32'hc1b820f3, 32'h4298aa17, 32'hc2bdf1e6};
test_label[798] = '{32'hc2049c76};
test_output[798] = '{32'h42daf8d4};
/*############ DEBUG ############
test_input[6384:6391] = '{18.2725727565, 29.9323834356, 17.4135187714, 69.41699268, -33.1527951686, -23.0160890596, 76.3322030039, -94.972454238};
test_label[798] = '{-33.1527951686};
test_output[798] = '{109.485990253};
############ END DEBUG ############*/
test_input[6392:6399] = '{32'h42b1dab3, 32'h41c4a5a2, 32'h42a0f7f2, 32'h429c82ac, 32'h427ad5ee, 32'h42a16e1f, 32'hc109be8e, 32'hc2c12644};
test_label[799] = '{32'h42b1dab3};
test_output[799] = '{32'h3a05a725};
/*############ DEBUG ############
test_input[6392:6399] = '{88.927143924, 24.5808758051, 80.48426621, 78.2552157814, 62.7089151721, 80.7150770929, -8.60902212049, -96.5747389052};
test_label[799] = '{88.927143924};
test_output[799] = '{0.000509845394713};
############ END DEBUG ############*/
test_input[6400:6407] = '{32'hc2611cdc, 32'h427d9db4, 32'hc2abc11c, 32'h42c72929, 32'hc25603ab, 32'hc2434f10, 32'h41e1b5a1, 32'h42b11dac};
test_label[800] = '{32'h42c72929};
test_output[800] = '{32'h3788fe95};
/*############ DEBUG ############
test_input[6400:6407] = '{-56.2781845605, 63.4040072379, -85.8771689616, 99.5803901902, -53.5035838887, -48.8272113132, 28.2136864564, 88.557953724};
test_label[800] = '{99.5803901902};
test_output[800] = '{1.63310128068e-05};
############ END DEBUG ############*/
test_input[6408:6415] = '{32'hc2b4e65c, 32'h41dcd5c4, 32'h424f3258, 32'hc1a587a7, 32'hbf6ccf8f, 32'hc280272d, 32'h41fe7774, 32'hc2c71b0e};
test_label[801] = '{32'hbf6ccf8f};
test_output[801] = '{32'h4252e596};
/*############ DEBUG ############
test_input[6408:6415] = '{-90.4499240386, 27.6043771731, 51.7991640306, -20.6912363955, -0.92504211041, -64.0765158044, 31.8083261865, -99.5528374627};
test_label[801] = '{-0.92504211041};
test_output[801] = '{52.7242061431};
############ END DEBUG ############*/
test_input[6416:6423] = '{32'hc2b8c311, 32'h411be96c, 32'hc2c3974e, 32'hc2707b40, 32'h42a1620f, 32'hc23bb2b7, 32'hc1119f08, 32'hc1a9b874};
test_label[802] = '{32'hc2707b40};
test_output[802] = '{32'h430ccfd8};
/*############ DEBUG ############
test_input[6416:6423] = '{-92.3809908308, 9.74448818452, -97.7955168219, -60.1203604515, 80.691522113, -46.9245253556, -9.10132620335, -21.215065425};
test_label[802] = '{-60.1203604515};
test_output[802] = '{140.811882565};
############ END DEBUG ############*/
test_input[6424:6431] = '{32'h427fd46a, 32'h41d5a04d, 32'h40085fc2, 32'hc2aa33c6, 32'h423ff641, 32'hbee6c210, 32'hc0ae24fc, 32'hc22d67c7};
test_label[803] = '{32'hc22d67c7};
test_output[803] = '{32'h42d69e18};
/*############ DEBUG ############
test_input[6424:6431] = '{63.9574362965, 26.7032723753, 2.13084449695, -85.1011231077, 47.9904820604, -0.45069932918, -5.44201482516, -43.3513435763};
test_label[803] = '{-43.3513435763};
test_output[803] = '{107.308779989};
############ END DEBUG ############*/
test_input[6432:6439] = '{32'h42a9eed7, 32'h42b034b4, 32'h425b6e1f, 32'hc2c06d43, 32'hc26d4dcc, 32'h4296f481, 32'hc2261ca9, 32'h422def8e};
test_label[804] = '{32'h422def8e};
test_output[804] = '{32'h4232a565};
/*############ DEBUG ############
test_input[6432:6439] = '{84.9664864932, 88.1029336695, 54.8575383358, -96.2134048924, -59.3259722967, 75.4775470442, -41.5279876618, 43.4839396878};
test_label[804] = '{43.4839396878};
test_output[804] = '{44.6615170582};
############ END DEBUG ############*/
test_input[6440:6447] = '{32'h42a5e34c, 32'h4056e0a5, 32'h429e2406, 32'h419dd4e6, 32'h41ac85fa, 32'h42b3cf1b, 32'hc252beac, 32'h4108ca16};
test_label[805] = '{32'h41ac85fa};
test_output[805] = '{32'h4288ae1b};
/*############ DEBUG ############
test_input[6440:6447] = '{82.943937884, 3.35746113827, 79.0703620332, 19.7289535664, 21.5654191351, 89.9045006154, -52.6862031404, 8.54933739288};
test_label[805] = '{21.5654191351};
test_output[805] = '{68.3400492893};
############ END DEBUG ############*/
test_input[6448:6455] = '{32'hc1ef5e41, 32'hc2a638f7, 32'hc18430c1, 32'h42af34f2, 32'hc2a77588, 32'h425639c0, 32'h4226e332, 32'hc299531a};
test_label[806] = '{32'h42af34f2};
test_output[806] = '{32'h26f00000};
/*############ DEBUG ############
test_input[6448:6455] = '{-29.9210223023, -83.1112569223, -16.5238057914, 87.6034087308, -83.72955083, 53.5563982229, 41.7218703102, -76.6623052527};
test_label[806] = '{87.6034087308};
test_output[806] = '{1.66533453694e-15};
############ END DEBUG ############*/
test_input[6456:6463] = '{32'h42529968, 32'h429f8483, 32'hc2707b3c, 32'hc1aa3ab6, 32'h422c2ea4, 32'hc26883b7, 32'hc26ef0ca, 32'hc27fabce};
test_label[807] = '{32'hc2707b3c};
test_output[807] = '{32'h430be110};
/*############ DEBUG ############
test_input[6456:6463] = '{52.6498117214, 79.7588116058, -60.1203454065, -21.2786681771, 43.0455490269, -58.1286261499, -59.7351469141, -63.917776262};
test_label[807] = '{-60.1203454065};
test_output[807] = '{139.879157012};
############ END DEBUG ############*/
test_input[6464:6471] = '{32'h42c25b00, 32'hc1cf4445, 32'hc12f2e31, 32'hc2769de5, 32'hc1fa5fc8, 32'hc21272e7, 32'h42afc4cb, 32'hc230a12f};
test_label[808] = '{32'hc1fa5fc8};
test_output[808] = '{32'h4300797f};
/*############ DEBUG ############
test_input[6464:6471] = '{97.1777368422, -25.9083339166, -10.948777377, -61.6541928335, -31.2967677552, -36.6122096518, 87.8843646449, -44.1574053402};
test_label[808] = '{-31.2967677552};
test_output[808] = '{128.474596625};
############ END DEBUG ############*/
test_input[6472:6479] = '{32'hc29d966b, 32'h4228d84f, 32'hc2b78bc1, 32'h42597fae, 32'hc1e8a17e, 32'hc27e154e, 32'hc0b2394d, 32'h4210c3e8};
test_label[809] = '{32'hc29d966b};
test_output[809] = '{32'h43052b21};
/*############ DEBUG ############
test_input[6472:6479] = '{-78.7937854274, 42.2112402966, -91.7729568921, 54.3746873863, -29.0788529154, -63.5208048169, -5.5694949206, 36.191313141};
test_label[809] = '{-78.7937854274};
test_output[809] = '{133.168478044};
############ END DEBUG ############*/
test_input[6480:6487] = '{32'hc25a7e67, 32'hc2b5dd11, 32'hc278cc4b, 32'h41480396, 32'h4271c078, 32'hc245dfa7, 32'hc2aa85ba, 32'hc2b14fe4};
test_label[810] = '{32'hc2aa85ba};
test_output[810] = '{32'h4311b2fb};
/*############ DEBUG ############
test_input[6480:6487] = '{-54.623440619, -90.9317687656, -62.1995046771, 12.5008758376, 60.43795768, -49.4684113267, -85.2611861559, -88.6560382258};
test_label[810] = '{-85.2611861559};
test_output[810] = '{145.699143836};
############ END DEBUG ############*/
test_input[6488:6495] = '{32'hc260b4a1, 32'h423bab02, 32'hc0dd6b06, 32'hc297e31a, 32'hc2ba2f44, 32'hc220b848, 32'h4274f74e, 32'hc2278770};
test_label[811] = '{32'hc2278770};
test_output[811] = '{32'h42ce3f5f};
/*############ DEBUG ############
test_input[6488:6495] = '{-56.1763955932, 46.9170016404, -6.91931420657, -75.9435546156, -93.0923189398, -40.1799610535, 61.2415072072, -41.8822629826};
test_label[811] = '{-41.8822629826};
test_output[811] = '{103.123770791};
############ END DEBUG ############*/
test_input[6496:6503] = '{32'hc134bd70, 32'hc1d36290, 32'hc2b071d4, 32'hc2263a50, 32'hc2af5dc4, 32'h42172e06, 32'hc29522e7, 32'h42561a1a};
test_label[812] = '{32'hc29522e7};
test_output[812] = '{32'h430017fa};
/*############ DEBUG ############
test_input[6496:6503] = '{-11.2962494294, -26.4231266557, -88.222317459, -41.5569448613, -87.683135989, 37.7949446469, -74.5681709428, 53.5254892273};
test_label[812] = '{-74.5681709428};
test_output[812] = '{128.093660317};
############ END DEBUG ############*/
test_input[6504:6511] = '{32'h41bd9465, 32'h42ae5775, 32'hc2ba1d8d, 32'h42019315, 32'h42603c08, 32'hc2baf340, 32'h418a7c07, 32'hc1f0872d};
test_label[813] = '{32'hc2ba1d8d};
test_output[813] = '{32'h43343a81};
/*############ DEBUG ############
test_input[6504:6511] = '{23.6974583807, 87.1708139402, -93.0577134157, 32.3936348226, 56.0586254897, -93.475100311, 17.3105604021, -30.0660037108};
test_label[813] = '{-93.0577134157};
test_output[813] = '{180.228527356};
############ END DEBUG ############*/
test_input[6512:6519] = '{32'h4230a06d, 32'h40c023c2, 32'hc2b24596, 32'hc26e798c, 32'hc2b357b7, 32'hc1d18055, 32'h42313b22, 32'hc1e68af7};
test_label[814] = '{32'h42313b22};
test_output[814] = '{32'h3f1ed64e};
/*############ DEBUG ############
test_input[6512:6519] = '{44.1566652809, 6.00436516239, -89.1359102434, -59.6186976753, -89.671315482, -26.187662684, 44.3077454124, -28.8178539206};
test_label[814] = '{44.3077454124};
test_output[814] = '{0.620457556192};
############ END DEBUG ############*/
test_input[6520:6527] = '{32'h41cebee1, 32'hc23c65c3, 32'hc1af741c, 32'h42880b72, 32'hc232e3f6, 32'hc2a85fa3, 32'hc21c8fea, 32'hc155dcbc};
test_label[815] = '{32'h41cebee1};
test_output[815] = '{32'h4228b774};
/*############ DEBUG ############
test_input[6520:6527] = '{25.843201766, -47.099377846, -21.9316934256, 68.0223566435, -44.7226181616, -84.1867921748, -39.1405404557, -13.3663898974};
test_label[815] = '{25.843201766};
test_output[815] = '{42.1791548775};
############ END DEBUG ############*/
test_input[6528:6535] = '{32'hc2a215dc, 32'h42347632, 32'h42ad7f0c, 32'h4228283e, 32'h42c31522, 32'hc226a206, 32'hc0bdb0b3, 32'h427ae6d1};
test_label[816] = '{32'h4228283e};
test_output[816] = '{32'h425e020b};
/*############ DEBUG ############
test_input[6528:6535] = '{-81.042694245, 45.1154269916, 86.7481420119, 42.0392987369, 97.5412747414, -41.6582272145, -5.92781969499, 62.7254067051};
test_label[816] = '{42.0392987369};
test_output[816] = '{55.5019965444};
############ END DEBUG ############*/
test_input[6536:6543] = '{32'h41a67e7a, 32'hc2a6b41d, 32'hc2693777, 32'h42c07926, 32'hc1412018, 32'hc26ffe55, 32'hc2538839, 32'hc065938c};
test_label[817] = '{32'h41a67e7a};
test_output[817] = '{32'h4296d987};
/*############ DEBUG ############
test_input[6536:6543] = '{20.8117560996, -83.3517850948, -58.3041652861, 96.236616595, -12.0703353008, -59.9983725629, -52.8830286264, -3.58713059642};
test_label[817] = '{20.8117560996};
test_output[817] = '{75.4248604954};
############ END DEBUG ############*/
test_input[6544:6551] = '{32'h42a58494, 32'h4218cce8, 32'h4287ab9f, 32'h42859cff, 32'hc1567bf9, 32'hc034d24d, 32'h41d1ef91, 32'hc2135832};
test_label[818] = '{32'h4218cce8};
test_output[818] = '{32'h42323c41};
/*############ DEBUG ############
test_input[6544:6551] = '{82.7589427018, 38.2001026625, 67.8351971816, 66.8066361254, -13.4052671554, -2.82533564357, 26.241976038, -36.8361267806};
test_label[818] = '{38.2001026625};
test_output[818] = '{44.5588404874};
############ END DEBUG ############*/
test_input[6552:6559] = '{32'hc25a71c4, 32'h428b0874, 32'h4137dc37, 32'h42016175, 32'hc1ccf9e7, 32'hc26bd6c3, 32'hc255e29a, 32'h411044e2};
test_label[819] = '{32'hc25a71c4};
test_output[819] = '{32'h42f84156};
/*############ DEBUG ############
test_input[6552:6559] = '{-54.6111011479, 69.5165114357, 11.4912632354, 32.3451722991, -25.6220224365, -58.9597282398, -53.4712913075, 9.01681744621};
test_label[819] = '{-54.6111011479};
test_output[819] = '{124.127612584};
############ END DEBUG ############*/
test_input[6560:6567] = '{32'hc2a7099f, 32'h41baa4dc, 32'h412064b6, 32'hc2176638, 32'h42c34042, 32'hc2868376, 32'h42722771, 32'h428d1baf};
test_label[820] = '{32'hc2176638};
test_output[820] = '{32'h430779af};
/*############ DEBUG ############
test_input[6560:6567] = '{-83.5187879261, 23.3304970646, 10.0245879499, -37.849824602, 97.6255049815, -67.2567588079, 60.5385166406, 70.5540692423};
test_label[820] = '{-37.849824602};
test_output[820] = '{135.475329584};
############ END DEBUG ############*/
test_input[6568:6575] = '{32'h42bbdea8, 32'hc213821e, 32'h42526837, 32'hc1a13120, 32'hc26de894, 32'h41a60d3c, 32'hc178c651, 32'h42627a6f};
test_label[821] = '{32'hc178c651};
test_output[821] = '{32'h42daf773};
/*############ DEBUG ############
test_input[6568:6575] = '{93.9348792687, -36.8770692338, 52.6017705162, -20.1489866553, -59.4771285798, 20.7564626851, -15.5484166937, 56.6195647381};
test_label[821] = '{-15.5484166937};
test_output[821] = '{109.483295962};
############ END DEBUG ############*/
test_input[6576:6583] = '{32'h4132941f, 32'h42a2ecb7, 32'h42095bbe, 32'h42bc322c, 32'hc247a130, 32'hc2c494a9, 32'hc29009b3, 32'hc0a1503b};
test_label[822] = '{32'hc0a1503b};
test_output[822] = '{32'h42c64730};
/*############ DEBUG ############
test_input[6576:6583] = '{11.1611627622, 81.4623341289, 34.3395922951, 94.0979889593, -49.9074098804, -98.2903483689, -72.0189407786, -5.04104381531};
test_label[822] = '{-5.04104381531};
test_output[822] = '{99.1390360285};
############ END DEBUG ############*/
test_input[6584:6591] = '{32'h427cb3f1, 32'hc172731d, 32'hc2afde3f, 32'h418a1a1e, 32'hc2816f6d, 32'hc212cf56, 32'hc2668d26, 32'h42a1b542};
test_label[823] = '{32'h427cb3f1};
test_output[823] = '{32'h418d6d27};
/*############ DEBUG ############
test_input[6584:6591] = '{63.1757224757, -15.1531034032, -87.9340721898, 17.2627519039, -64.7176313281, -36.702478018, -57.6378389356, 80.8540192704};
test_label[823] = '{63.1757224757};
test_output[823] = '{17.6782968157};
############ END DEBUG ############*/
test_input[6592:6599] = '{32'hc2bd43ad, 32'hc251cfd3, 32'h4218699f, 32'hc23c2a69, 32'h409ba4e8, 32'hc22798b6, 32'h3e5d7a81, 32'hc22c52c0};
test_label[824] = '{32'h3e5d7a81};
test_output[824] = '{32'h42178c24};
/*############ DEBUG ############
test_input[6592:6599] = '{-94.6321810153, -52.4529521373, 38.1031439391, -47.0414156676, 4.8638801946, -41.8991310078, 0.21628763289, -43.0808089662};
test_label[824] = '{0.21628763289};
test_output[824] = '{37.8868563062};
############ END DEBUG ############*/
test_input[6600:6607] = '{32'hc189be7a, 32'h400205c8, 32'hc217bd3b, 32'h42abd835, 32'hc262f774, 32'h42a86d40, 32'h42071abb, 32'hc2487921};
test_label[825] = '{32'hc2487921};
test_output[825] = '{32'h430834fd};
/*############ DEBUG ############
test_input[6600:6607] = '{-17.2180062908, 2.03160280983, -37.9347953637, 85.9222777825, -56.7416540647, 84.2133810305, 33.7761044417, -50.1182882471};
test_label[825] = '{-50.1182882471};
test_output[825] = '{136.206982978};
############ END DEBUG ############*/
test_input[6608:6615] = '{32'hc2020c29, 32'h428559c3, 32'h41aa8fb8, 32'hc2a590e5, 32'h42b52b3a, 32'h42599fa9, 32'hc1081553, 32'h41ca4fe4};
test_label[826] = '{32'h41ca4fe4};
test_output[826] = '{32'h42829741};
/*############ DEBUG ############
test_input[6608:6615] = '{-32.5118743854, 66.6753130496, 21.3201750152, -82.7829984483, 90.5844300784, 54.4059192428, -8.50520603034, 25.2890090759};
test_label[826] = '{25.2890090759};
test_output[826] = '{65.2954210025};
############ END DEBUG ############*/
test_input[6616:6623] = '{32'hc2660508, 32'hc2be3451, 32'hc26c69a1, 32'h428d2dfd, 32'h41e6a7c1, 32'h42a04681, 32'h415cd4ac, 32'h4181305a};
test_label[827] = '{32'hc26c69a1};
test_output[827] = '{32'h430b3dae};
/*############ DEBUG ############
test_input[6616:6623] = '{-57.5049142464, -95.1021799349, -59.103153371, 70.5898199955, 28.8319117558, 80.1377047366, 13.8019217801, 16.1486084874};
test_label[827] = '{-59.103153371};
test_output[827] = '{139.240929457};
############ END DEBUG ############*/
test_input[6624:6631] = '{32'hc29890e7, 32'hc227ba66, 32'hc277e02f, 32'hc29f74ee, 32'hc29b48ae, 32'h423846da, 32'h4266d87f, 32'hc1a065be};
test_label[828] = '{32'h4266d87f};
test_output[828] = '{32'h37136c0e};
/*############ DEBUG ############
test_input[6624:6631] = '{-76.2830130919, -41.9320299035, -61.9689291684, -79.728376225, -77.6419522448, 46.0691924197, 57.7114205623, -20.0496780708};
test_label[828] = '{57.7114205623};
test_output[828] = '{8.78704099386e-06};
############ END DEBUG ############*/
test_input[6632:6639] = '{32'h41e85797, 32'hc2bc4883, 32'hc2349a90, 32'hc1b532bb, 32'hc2987188, 32'hc2c3eccd, 32'hc245a38d, 32'hc29de4e0};
test_label[829] = '{32'hc2349a90};
test_output[829] = '{32'h4294632e};
/*############ DEBUG ############
test_input[6632:6639] = '{29.0427690859, -94.1416220991, -45.1509406987, -22.6497708075, -76.2217410689, -97.9624994854, -49.4097181458, -78.9470179721};
test_label[829] = '{-45.1509406987};
test_output[829] = '{74.1937097846};
############ END DEBUG ############*/
test_input[6640:6647] = '{32'h428147a6, 32'hc0f262d7, 32'h42b7bccc, 32'h42796cd5, 32'hc20b1464, 32'hc19a2a07, 32'h429fcf5b, 32'hc27852ad};
test_label[830] = '{32'hc20b1464};
test_output[830] = '{32'h42fd46ff};
/*############ DEBUG ############
test_input[6640:6647] = '{64.6399411092, -7.57456550171, 91.8687474909, 62.3562819948, -34.769913581, -19.2705215598, 79.9049910728, -62.0807396033};
test_label[830] = '{-34.769913581};
test_output[830] = '{126.638667443};
############ END DEBUG ############*/
test_input[6648:6655] = '{32'h42a96aac, 32'h428f7719, 32'hc2af81a6, 32'hc2b8be3a, 32'h4226ead1, 32'h420ea94b, 32'hc264fc97, 32'h42996aa2};
test_label[831] = '{32'h420ea94b};
test_output[831] = '{32'h42442c66};
/*############ DEBUG ############
test_input[6648:6655] = '{84.7083458108, 71.7326145901, -87.7532225802, -92.3715395383, 41.7293116974, 35.6653269355, -57.2466701623, 76.7082636586};
test_label[831] = '{35.6653269355};
test_output[831] = '{49.0433565692};
############ END DEBUG ############*/
test_input[6656:6663] = '{32'h429b19aa, 32'h41708a26, 32'hc2472ec3, 32'hc286dd23, 32'h4235f018, 32'h42a711fb, 32'h42aee922, 32'hc28cdf7d};
test_label[832] = '{32'hc286dd23};
test_output[832] = '{32'h431ae82d};
/*############ DEBUG ############
test_input[6656:6663] = '{77.5501236531, 15.0337275197, -49.7956661827, -67.4319042716, 45.4844681639, 83.5351142886, 87.4553364377, -70.4364974095};
test_label[832] = '{-67.4319042716};
test_output[832] = '{154.906932155};
############ END DEBUG ############*/
test_input[6664:6671] = '{32'h41eb8469, 32'hc23fd9af, 32'h422cd30b, 32'h423982be, 32'h41905623, 32'h42a67898, 32'h429f5343, 32'h42a1b803};
test_label[833] = '{32'h429f5343};
test_output[833] = '{32'h406bf9c2};
/*############ DEBUG ############
test_input[6664:6671] = '{29.4396541453, -47.9625824707, 43.2060983628, 46.3776788869, 18.042059664, 83.2355370656, 79.6626235321, 80.8593976912};
test_label[833] = '{79.6626235321};
test_output[833] = '{3.68711907645};
############ END DEBUG ############*/
test_input[6672:6679] = '{32'hc19c69d9, 32'hc28f1426, 32'hc2b9303c, 32'hc1486199, 32'hbf569af6, 32'hc2450f29, 32'hc2a6eb34, 32'h410b4439};
test_label[834] = '{32'hc1486199};
test_output[834] = '{32'h41a9d30e};
/*############ DEBUG ############
test_input[6672:6679] = '{-19.5516843686, -71.5393490166, -92.5942044819, -12.5238273637, -0.83830200703, -49.2648063318, -83.4593803192, 8.70415575915};
test_label[834] = '{-12.5238273637};
test_output[834] = '{21.2280548611};
############ END DEBUG ############*/
test_input[6680:6687] = '{32'hc2747f76, 32'hc2b7a16a, 32'hc2bc855a, 32'h42a337ef, 32'h422733c0, 32'h422d3437, 32'hc20ff182, 32'h42aae927};
test_label[835] = '{32'hc2747f76};
test_output[835] = '{32'h431299db};
/*############ DEBUG ############
test_input[6680:6687] = '{-61.1244743862, -91.8152650448, -94.2604527973, 81.6092455428, 41.8005353009, 43.3009901823, -35.9858462875, 85.4553790572};
test_label[835] = '{-61.1244743862};
test_output[835] = '{146.600990644};
############ END DEBUG ############*/
test_input[6688:6695] = '{32'h42af0c04, 32'h4218ea93, 32'h426eaf79, 32'h41eb7006, 32'hc2b47780, 32'h4180d8c2, 32'h4298b5e1, 32'h42ad7057};
test_label[836] = '{32'hc2b47780};
test_output[836] = '{32'h43322071};
/*############ DEBUG ############
test_input[6688:6695] = '{87.5234714352, 38.2290762821, 59.6713612868, 29.4296994627, -90.2333998644, 16.1058395719, 76.3552328269, 86.7194122105};
test_label[836] = '{-90.2333998644};
test_output[836] = '{178.126725015};
############ END DEBUG ############*/
test_input[6696:6703] = '{32'hc0400fcf, 32'h41fe3f73, 32'h422fe0cf, 32'h412bb24c, 32'h418aa4ab, 32'hc29690a9, 32'hc202734e, 32'hc1ee1da0};
test_label[837] = '{32'h412bb24c};
test_output[837] = '{32'h4204f43e};
/*############ DEBUG ############
test_input[6696:6703] = '{-3.00096479297, 31.7809802382, 43.9695406799, 10.7310297517, 17.3304039249, -75.282542341, -32.6126012792, -29.7644649316};
test_label[837] = '{10.7310297517};
test_output[837] = '{33.2385160166};
############ END DEBUG ############*/
test_input[6704:6711] = '{32'h421aae8a, 32'h418c6803, 32'h42c1cc84, 32'hc2acc40e, 32'h42a6f4cf, 32'h418e0d6c, 32'h418aef5d, 32'hc29fa2c1};
test_label[838] = '{32'h42c1cc84};
test_output[838] = '{32'h35c7128c};
/*############ DEBUG ############
test_input[6704:6711] = '{38.6704480666, 17.5507871753, 96.8994471623, -86.3829176042, 83.4781428446, 17.7565541507, 17.36687636, -79.8178798605};
test_label[838] = '{96.8994471623};
test_output[838] = '{1.48320531406e-06};
############ END DEBUG ############*/
test_input[6712:6719] = '{32'h42a1e620, 32'hc1a928d7, 32'hc2a8c329, 32'h425158d9, 32'hc225eea1, 32'hc190230c, 32'hc12ae8f3, 32'hc275df78};
test_label[839] = '{32'hc225eea1};
test_output[839] = '{32'h42f4dd71};
/*############ DEBUG ############
test_input[6712:6719] = '{80.9494646869, -21.144941392, -84.3811684111, 52.3367643854, -41.4830357781, -18.0171129711, -10.6818724382, -61.4682299467};
test_label[839] = '{-41.4830357781};
test_output[839] = '{122.432500465};
############ END DEBUG ############*/
test_input[6720:6727] = '{32'h42c014c8, 32'hc1e1599b, 32'hc1b04587, 32'h3fa6ad3c, 32'h41ac1d55, 32'h429c2c85, 32'h427780ff, 32'h41346086};
test_label[840] = '{32'h42c014c8};
test_output[840] = '{32'h32890855};
/*############ DEBUG ############
test_input[6720:6727] = '{96.0405879359, -28.1687529194, -22.0339491753, 1.30216173579, 21.5143214437, 78.0869493096, 61.8759711992, 11.2735650015};
test_label[840] = '{96.0405879359};
test_output[840] = '{1.59526871875e-08};
############ END DEBUG ############*/
test_input[6728:6735] = '{32'hc2482a14, 32'hc232bf73, 32'hc2a00206, 32'h401fbe54, 32'hc20a28d0, 32'h4299b508, 32'hc09a8560, 32'hc1f3e32a};
test_label[841] = '{32'hc20a28d0};
test_output[841] = '{32'h42dec970};
/*############ DEBUG ############
test_input[6728:6735] = '{-50.041091153, -44.6869627977, -80.0039544682, 2.49599163622, -34.539855487, 76.8535797056, -4.82878116209, -30.4859201603};
test_label[841] = '{-34.539855487};
test_output[841] = '{111.393435193};
############ END DEBUG ############*/
test_input[6736:6743] = '{32'hc11d59e0, 32'h4287f182, 32'hc2bca337, 32'h4287e214, 32'hc1bbf7a1, 32'h429616ea, 32'h42b26506, 32'h4229db98};
test_label[842] = '{32'hc1bbf7a1};
test_output[842] = '{32'h42e162ef};
/*############ DEBUG ############
test_input[6736:6743] = '{-9.83444174266, 67.9716927442, -94.3187760995, 67.941561465, -23.4959117736, 75.0447508596, 89.1973142182, 42.4644485972};
test_label[842] = '{-23.4959117736};
test_output[842] = '{112.693226707};
############ END DEBUG ############*/
test_input[6744:6751] = '{32'h426867ac, 32'hc2673ca7, 32'h42bbd2bd, 32'h41d308c8, 32'hc1d0eaed, 32'hc2bf70aa, 32'hc20dffbc, 32'hc1bf9b98};
test_label[843] = '{32'hc2bf70aa};
test_output[843] = '{32'h433da1b4};
/*############ DEBUG ############
test_input[6744:6751] = '{58.1012422529, -57.8092327111, 93.9115957952, 26.3792871174, -26.1147089591, -95.7200494296, -35.4997420828, -23.9509733903};
test_label[843] = '{-95.7200494296};
test_output[843] = '{189.631645225};
############ END DEBUG ############*/
test_input[6752:6759] = '{32'hc257d562, 32'h41c5d024, 32'hc299b4bd, 32'hc1cd7df6, 32'h4179dec4, 32'hc2905eb0, 32'hc253e751, 32'hc2969878};
test_label[844] = '{32'h4179dec4};
test_output[844] = '{32'h4111c1f8};
/*############ DEBUG ############
test_input[6752:6759] = '{-53.9583807254, 24.7266311764, -76.8530054076, -25.6865036925, 15.6168865103, -72.1849379257, -52.9758943183, -75.297787754};
test_label[844] = '{15.6168865103};
test_output[844] = '{9.10985524298};
############ END DEBUG ############*/
test_input[6760:6767] = '{32'hc2b01797, 32'h418924a8, 32'hc0a574dd, 32'h425817ef, 32'h414c129f, 32'h42775024, 32'h42a28131, 32'hc20e2cc1};
test_label[845] = '{32'h414c129f};
test_output[845] = '{32'h4288fedd};
/*############ DEBUG ############
test_input[6760:6767] = '{-88.0460709049, 17.1428977003, -5.17051571998, 54.0233709735, 12.7545464912, 61.8282640634, 81.2523254038, -35.54370639};
test_label[845] = '{12.7545464912};
test_output[845] = '{68.4977789162};
############ END DEBUG ############*/
test_input[6768:6775] = '{32'hc225b885, 32'h429af0f3, 32'hc2b05404, 32'h4132266d, 32'hc29a99cd, 32'h42c3ba73, 32'h42002332, 32'h423521fd};
test_label[846] = '{32'hc225b885};
test_output[846] = '{32'h430b4b5b};
/*############ DEBUG ############
test_input[6768:6775] = '{-41.4301936997, 77.4706054286, -88.1640964477, 11.1343816711, -77.3003886356, 97.864160956, 32.0343713885, 45.2831934598};
test_label[846] = '{-41.4301936997};
test_output[846] = '{139.294354657};
############ END DEBUG ############*/
test_input[6776:6783] = '{32'h41c97f9d, 32'h42c269f5, 32'h413b5614, 32'h42c3d807, 32'hc2820c8a, 32'h4258018d, 32'h4108bdca, 32'hc23010f1};
test_label[847] = '{32'h4258018d};
test_output[847] = '{32'h4231464d};
/*############ DEBUG ############
test_input[6776:6783] = '{25.1873117139, 97.2069450848, 11.7085148331, 97.9219321768, -65.0244895127, 54.0015162014, 8.54633555977, -44.0165437532};
test_label[847] = '{54.0015162014};
test_output[847] = '{44.3186539817};
############ END DEBUG ############*/
test_input[6784:6791] = '{32'h42352237, 32'hc202945b, 32'hc223868d, 32'hc2c775c3, 32'hc2273def, 32'hc24987d8, 32'h4215f807, 32'h428b293a};
test_label[848] = '{32'hc223868d};
test_output[848] = '{32'h42dcec80};
/*############ DEBUG ############
test_input[6784:6791] = '{45.2834117436, -32.6448797757, -40.8813966183, -99.7300005129, -41.8104813256, -50.382659258, 37.4922142992, 69.5805192077};
test_label[848] = '{-40.8813966183};
test_output[848] = '{110.461915826};
############ END DEBUG ############*/
test_input[6792:6799] = '{32'h41e3bca1, 32'hc23a1810, 32'h4161217e, 32'h415462bd, 32'hc29b8eac, 32'h425b1d77, 32'hc20d7f4d, 32'h4290add0};
test_label[849] = '{32'h425b1d77};
test_output[849] = '{32'h418c7c52};
/*############ DEBUG ############
test_input[6792:6799] = '{28.4671047817, -46.5234978904, 14.0706764899, 13.2741058543, -77.7786550517, 54.778774847, -35.3743179908, 72.3394785033};
test_label[849] = '{54.778774847};
test_output[849] = '{17.56070368};
############ END DEBUG ############*/
test_input[6800:6807] = '{32'h42021d05, 32'hc2375231, 32'hc2c3fe96, 32'h42563337, 32'h4263c304, 32'h4223a4fa, 32'hc2c743cd, 32'h426e8d81};
test_label[850] = '{32'hc2c3fe96};
test_output[850] = '{32'h431db3e7};
/*############ DEBUG ############
test_input[6800:6807] = '{32.5283409079, -45.830266492, -97.9972389141, 53.5500159933, 56.9404432462, 40.9111089421, -99.6324244359, 59.6381888777};
test_label[850] = '{-97.9972389141};
test_output[850] = '{157.702737547};
############ END DEBUG ############*/
test_input[6808:6815] = '{32'hc29a3a12, 32'h42ba227c, 32'hc1dce44d, 32'hc2138388, 32'h42a196e4, 32'hbf008e5c, 32'h423016d1, 32'h4283aa08};
test_label[851] = '{32'h42ba227c};
test_output[851] = '{32'h369cf74c};
/*############ DEBUG ############
test_input[6808:6815] = '{-77.1134177037, 93.0673556818, -27.6114758279, -36.8784490755, 80.7947074354, -0.502172225864, 44.0222812198, 65.8320948887};
test_label[851] = '{93.0673556818};
test_output[851] = '{4.67795145189e-06};
############ END DEBUG ############*/
test_input[6816:6823] = '{32'h3e51f443, 32'hc291a877, 32'h4283ebec, 32'hc2762621, 32'h40d56670, 32'h417384ad, 32'h42874cdc, 32'hc1ed3238};
test_label[852] = '{32'h42874cdc};
test_output[852] = '{32'h3e2d823f};
/*############ DEBUG ############
test_input[6816:6823] = '{0.205033349998, -72.8290345072, 65.960788167, -61.5372368152, 6.66875471561, 15.2198911477, 67.6501147392, -29.6495207936};
test_label[852] = '{67.6501147392};
test_output[852] = '{0.169442160993};
############ END DEBUG ############*/
test_input[6824:6831] = '{32'h41d3635d, 32'hc11f3f28, 32'hc2ab2dbc, 32'h4293f4f8, 32'h4217fbc0, 32'hc25bbebc, 32'hc2a8be98, 32'h42819890};
test_label[853] = '{32'hc11f3f28};
test_output[853] = '{32'h42a7dceb};
/*############ DEBUG ############
test_input[6824:6831] = '{26.42351705, -9.95291922154, -85.5893249029, 73.9784572284, 37.9958493517, -54.9362655965, -84.3722533174, 64.7979733101};
test_label[853] = '{-9.95291922154};
test_output[853] = '{83.9314794753};
############ END DEBUG ############*/
test_input[6832:6839] = '{32'hc2b0d528, 32'hc2a5f891, 32'hc1a7bc0d, 32'h3f54cc85, 32'hc09fc127, 32'h41c97dd5, 32'h42c7842f, 32'hc2a06829};
test_label[854] = '{32'hc2b0d528};
test_output[854] = '{32'h433c2cac};
/*############ DEBUG ############
test_input[6832:6839] = '{-88.4163240035, -82.9854810383, -20.9668219481, 0.83124571917, -4.99232817311, 25.1864409597, 99.7581700134, -80.2034404645};
test_label[854] = '{-88.4163240035};
test_output[854] = '{188.174494017};
############ END DEBUG ############*/
test_input[6840:6847] = '{32'hc1832f97, 32'hc0c757bf, 32'h423cf181, 32'hc2878d76, 32'h428b4775, 32'h410f97cd, 32'hc1aa9e74, 32'hc1af5903};
test_label[855] = '{32'hc1832f97};
test_output[855] = '{32'h42ac135b};
/*############ DEBUG ############
test_input[6840:6847] = '{-16.3982365329, -6.22946119692, 47.2358424857, -67.7762923812, 69.6395676804, 8.97456073528, -21.3273698337, -21.9184625846};
test_label[855] = '{-16.3982365329};
test_output[855] = '{86.0378042135};
############ END DEBUG ############*/
test_input[6848:6855] = '{32'hc16c58aa, 32'hc2173f08, 32'hc236a686, 32'h41596131, 32'h423adccb, 32'h4285506f, 32'hc280c47c, 32'h421e8ca2};
test_label[856] = '{32'h421e8ca2};
test_output[856] = '{32'h41d8287a};
/*############ DEBUG ############
test_input[6848:6855] = '{-14.7716464569, -37.8115533959, -45.6626194164, 13.5862281467, 46.7156166316, 66.6570998066, -64.3837615247, 39.6373357163};
test_label[856] = '{39.6373357163};
test_output[856] = '{27.0197640925};
############ END DEBUG ############*/
test_input[6856:6863] = '{32'hc2a68853, 32'hc1e12028, 32'h426970fb, 32'hc28ab1f2, 32'h424a19b8, 32'hc26c15a4, 32'h4215d8dd, 32'h42b97e30};
test_label[857] = '{32'hc26c15a4};
test_output[857] = '{32'h4317c481};
/*############ DEBUG ############
test_input[6856:6863] = '{-83.2662570374, -28.1407017641, 58.3603308623, -69.347551272, 50.5251144407, -59.0211316042, 37.4617806857, 92.7464612759};
test_label[857] = '{-59.0211316042};
test_output[857] = '{151.76759288};
############ END DEBUG ############*/
test_input[6864:6871] = '{32'hc19d9124, 32'hc20de93e, 32'hc252045a, 32'hc170464d, 32'h4256fc9d, 32'hc27aab92, 32'hc171e0a4, 32'hc20dacd2};
test_label[858] = '{32'hc171e0a4};
test_output[858] = '{32'h4289ba63};
/*############ DEBUG ############
test_input[6864:6871] = '{-19.6958700789, -35.4777743765, -52.5042491036, -15.0171633884, 53.746694443, -62.6675473483, -15.1173440702, -35.4187690271};
test_label[858] = '{-15.1173440702};
test_output[858] = '{68.8640385133};
############ END DEBUG ############*/
test_input[6872:6879] = '{32'h42048c09, 32'hc29d00a9, 32'h42b4a981, 32'hc281a674, 32'hc114e83f, 32'h42a6a95b, 32'hc289668f, 32'hc24f4fd1};
test_label[859] = '{32'hc29d00a9};
test_output[859] = '{32'h4328d551};
/*############ DEBUG ############
test_input[6872:6879] = '{33.1367516519, -78.5012919673, 90.3310616201, -64.8251049101, -9.30670113154, 83.3307747428, -68.7003111097, -51.8279474151};
test_label[859] = '{-78.5012919673};
test_output[859] = '{168.833264793};
############ END DEBUG ############*/
test_input[6880:6887] = '{32'hc23d294b, 32'hc1cdf357, 32'hc28bc922, 32'hc2b88221, 32'h41386418, 32'hc2515a9e, 32'h4261de2f, 32'h42287bda};
test_label[860] = '{32'hc28bc922};
test_output[860] = '{32'h42fcb83a};
/*############ DEBUG ############
test_input[6880:6887] = '{-47.2903254706, -25.7438183148, -69.8928408861, -92.2541603238, 11.5244366896, -52.3384945204, 56.4669754357, 42.1209482341};
test_label[860] = '{-69.8928408861};
test_output[860] = '{126.35981691};
############ END DEBUG ############*/
test_input[6888:6895] = '{32'h429cce5e, 32'h429f6329, 32'h406a93cd, 32'h423ac9e2, 32'hc2b0f549, 32'h41019089, 32'h42832373, 32'h41cf4665};
test_label[861] = '{32'h41cf4665};
test_output[861] = '{32'h42581bfb};
/*############ DEBUG ############
test_input[6888:6895] = '{78.4030589359, 79.6936689982, 3.66527106535, 46.697150298, -88.4790743671, 8.09778709656, 65.5692393419, 25.9093732706};
test_label[861] = '{25.9093732706};
test_output[861] = '{54.0273231863};
############ END DEBUG ############*/
test_input[6896:6903] = '{32'h429aa1db, 32'hc2aa5300, 32'hc2bd785d, 32'hc285eaff, 32'hc16b551b, 32'h429823a8, 32'h427aa8f3, 32'hc2ba0b64};
test_label[862] = '{32'hc2aa5300};
test_output[862] = '{32'h4322bb1f};
/*############ DEBUG ############
test_input[6896:6903] = '{77.3161262822, -85.1621075896, -94.7350839329, -66.9589756493, -14.708277908, 76.0696439169, 62.6649899866, -93.0222501223};
test_label[862] = '{-85.1621075896};
test_output[862] = '{162.730947739};
############ END DEBUG ############*/
test_input[6904:6911] = '{32'hc2108dbd, 32'h42a7cf2a, 32'h4291970a, 32'h426b89b9, 32'h425b6792, 32'h41f1cebb, 32'h40da46f3, 32'hc2a038fa};
test_label[863] = '{32'h4291970a};
test_output[863] = '{32'h4131c117};
/*############ DEBUG ############
test_input[6904:6911] = '{-36.138417841, 83.9046210743, 72.7949953848, 58.8844932329, 54.8511434021, 30.2259428448, 6.82116078644, -80.1112841024};
test_label[863] = '{72.7949953848};
test_output[863] = '{11.109640657};
############ END DEBUG ############*/
test_input[6912:6919] = '{32'h4188297d, 32'hc28213d4, 32'h41bf19e4, 32'hc27997dc, 32'h3fd2b6ae, 32'h42a3b420, 32'h42b1ff29, 32'hc2b998b6};
test_label[864] = '{32'h42a3b420};
test_output[864] = '{32'h40e4b6f4};
/*############ DEBUG ############
test_input[6912:6919] = '{17.0202570687, -65.0387246871, 23.8876417752, -62.3983020613, 1.64619997328, 81.8518102998, 88.9983559392, -92.7982641446};
test_label[864] = '{81.8518102998};
test_output[864] = '{7.14733290933};
############ END DEBUG ############*/
test_input[6920:6927] = '{32'hc1a08972, 32'hc2b3004f, 32'hc268ef8f, 32'h426f9809, 32'h4211a312, 32'hc2b0985b, 32'h422750c0, 32'hc13066fa};
test_label[865] = '{32'hc2b0985b};
test_output[865] = '{32'h43143230};
/*############ DEBUG ############
test_input[6920:6927] = '{-20.0671121542, -89.5006034213, -58.2339430895, 59.8984725683, 36.4092480768, -88.2975691788, 41.8288581105, -11.0251409177};
test_label[865] = '{-88.2975691788};
test_output[865] = '{148.196041761};
############ END DEBUG ############*/
test_input[6928:6935] = '{32'h42a56c0f, 32'hbf04240f, 32'h422dd0be, 32'h423675ea, 32'h42b38f17, 32'h42c62ed5, 32'h427fb3b6, 32'h4289ff15};
test_label[866] = '{32'h423675ea};
test_output[866] = '{32'h4255e7d9};
/*############ DEBUG ############
test_input[6928:6935] = '{82.7110548083, -0.516175191387, 43.4538493708, 45.6151497204, 89.7794746882, 99.0914718192, 63.9254978688, 68.9982103234};
test_label[866] = '{45.6151497204};
test_output[866] = '{53.4764125055};
############ END DEBUG ############*/
test_input[6936:6943] = '{32'h4290977d, 32'hc2958f9a, 32'hc29e1dd2, 32'h40c905fc, 32'hc204cd47, 32'hc20cfb46, 32'hc290df93, 32'hc2bd3ded};
test_label[867] = '{32'hc2bd3ded};
test_output[867] = '{32'h4326eab5};
/*############ DEBUG ############
test_input[6936:6943] = '{72.2958722444, -74.7804720353, -79.0582450547, 6.28198040325, -33.200466252, -35.245385218, -72.4366687818, -94.6209501422};
test_label[867] = '{-94.6209501422};
test_output[867] = '{166.916822387};
############ END DEBUG ############*/
test_input[6944:6951] = '{32'hc2b8ac29, 32'hc148109f, 32'h42951cee, 32'h42c2037f, 32'hc2b1bf6d, 32'hc233faca, 32'hc29a3f60, 32'h425c713b};
test_label[868] = '{32'hc29a3f60};
test_output[868] = '{32'h432e216f};
/*############ DEBUG ############
test_input[6944:6951] = '{-92.3362527286, -12.5040577981, 74.5565020806, 97.0068262711, -88.8738790018, -44.9949130002, -77.1237792723, 55.1105753092};
test_label[868] = '{-77.1237792723};
test_output[868] = '{174.130605544};
############ END DEBUG ############*/
test_input[6952:6959] = '{32'hc08b852c, 32'hc2477ad1, 32'hc24528a9, 32'hc006cd8a, 32'hc2bfe3c6, 32'hc04a35c3, 32'hc1cb0ca1, 32'h40390828};
test_label[869] = '{32'h40390828};
test_output[869] = '{32'h3c201f8c};
/*############ DEBUG ############
test_input[6952:6959] = '{-4.36000616325, -49.869938133, -49.2897073801, -2.106295195, -95.9448704465, -3.15953131122, -25.3811667815, 2.89112285068};
test_label[869] = '{2.89112285068};
test_output[869] = '{0.00977314652468};
############ END DEBUG ############*/
test_input[6960:6967] = '{32'hc29363ec, 32'hc0762071, 32'h4272f1e5, 32'h41cf8987, 32'hc2982145, 32'h42893918, 32'h429dd865, 32'h4212ab3f};
test_label[870] = '{32'h4272f1e5};
test_output[870] = '{32'h41917ddb};
/*############ DEBUG ############
test_input[6960:6967] = '{-73.6951575187, -3.84572999633, 60.7362244612, 25.9421515482, -76.0649822906, 68.6115094798, 78.9226433946, 36.667233919};
test_label[870] = '{60.7362244612};
test_output[870] = '{18.1864522061};
############ END DEBUG ############*/
test_input[6968:6975] = '{32'h4099e933, 32'hc24c5360, 32'hc21f1032, 32'hc12c42ea, 32'hc2329006, 32'h4295d7f7, 32'h42983489, 32'hc201c6da};
test_label[871] = '{32'h42983489};
test_output[871] = '{32'h3e8917c9};
/*############ DEBUG ############
test_input[6968:6975] = '{4.80971669346, -51.0814227067, -39.7658147862, -10.7663366754, -44.6406497203, 74.9218073042, 76.1026077821, -32.4441894007};
test_label[871] = '{76.1026077821};
test_output[871] = '{0.267759581367};
############ END DEBUG ############*/
test_input[6976:6983] = '{32'hc22e1e98, 32'h4219df46, 32'h42aecf31, 32'hc1ae59a6, 32'hc25d91a9, 32'h42bb902d, 32'hc1339127, 32'hc27ec7ab};
test_label[872] = '{32'h4219df46};
test_output[872] = '{32'h425d42d1};
/*############ DEBUG ############
test_input[6976:6983] = '{-43.5298770519, 38.468039411, 87.4046692282, -21.7937741843, -55.3922478986, 93.7815910965, -11.2229379941, -63.6949883258};
test_label[872] = '{38.468039411};
test_output[872] = '{55.3152505904};
############ END DEBUG ############*/
test_input[6984:6991] = '{32'h424408c7, 32'h41facea0, 32'h42834f9b, 32'h41fb661a, 32'h42a1d644, 32'hc2112512, 32'h40dedf24, 32'hbf18e5d5};
test_label[873] = '{32'h424408c7};
test_output[873] = '{32'h41ff4781};
/*############ DEBUG ############
test_input[6984:6991] = '{49.0085729751, 31.350891497, 65.6554758538, 31.4248543161, 80.9184868499, -36.2862024657, 6.96473866916, -0.597256987038};
test_label[873] = '{49.0085729751};
test_output[873] = '{31.90991411};
############ END DEBUG ############*/
test_input[6992:6999] = '{32'hc2aa1ea2, 32'h415c6bf1, 32'hc1c20d48, 32'hbf45f898, 32'hc2b8ca80, 32'h411c3567, 32'hc292475f, 32'hc0d10839};
test_label[874] = '{32'hc2aa1ea2};
test_output[874] = '{32'h42c5b54c};
/*############ DEBUG ############
test_input[6992:6999] = '{-85.0598323945, 13.7763530808, -24.2564852646, -0.77332449531, -92.3955083816, 9.76303738726, -73.1393938512, -6.53225386503};
test_label[874] = '{-85.0598323945};
test_output[874] = '{98.8540979364};
############ END DEBUG ############*/
test_input[7000:7007] = '{32'hc2b0ba6a, 32'hc1dde6e2, 32'h4272563e, 32'h41f06ba2, 32'hc26b3976, 32'hc255c285, 32'h42a5a216, 32'hc21b49da};
test_label[875] = '{32'h4272563e};
test_output[875] = '{32'h41b1dbdd};
/*############ DEBUG ############
test_input[7000:7007] = '{-88.3640918218, -27.7377364845, 60.5842201182, 30.0525542387, -58.8061157717, -53.4399588582, 82.8165748551, -38.8221196773};
test_label[875] = '{60.5842201182};
test_output[875] = '{22.2323547371};
############ END DEBUG ############*/
test_input[7008:7015] = '{32'hc2579b79, 32'hc2352a4f, 32'hc29d5786, 32'h42616921, 32'hc228ab4a, 32'hc2b2828a, 32'hc1c39043, 32'hc18b7df5};
test_label[876] = '{32'hc1c39043};
test_output[876] = '{32'h42a198a1};
/*############ DEBUG ############
test_input[7008:7015] = '{-53.901830087, -45.2913187636, -78.6709445846, 56.3526654535, -42.1672740782, -89.2549614689, -24.4454400786, -17.4365029915};
test_label[876] = '{-24.4454400786};
test_output[876] = '{80.7981055321};
############ END DEBUG ############*/
test_input[7016:7023] = '{32'hc2b7b2f9, 32'h421f0524, 32'h3fdf3e60, 32'h4284cc51, 32'h41e1b640, 32'h408d53f1, 32'h4259bb49, 32'h424a9d22};
test_label[877] = '{32'h4259bb49};
test_output[877] = '{32'h413f7569};
/*############ DEBUG ############
test_input[7016:7023] = '{-91.8495549763, 39.7550186762, 1.74409099575, 66.3990528704, 28.2139894485, 4.41649689287, 54.4328949735, 50.6534502596};
test_label[877] = '{54.4328949735};
test_output[877] = '{11.9661643977};
############ END DEBUG ############*/
test_input[7024:7031] = '{32'hc28f9faa, 32'hc2504d51, 32'hc0ece64f, 32'h4242be9d, 32'h4187a01b, 32'h41253406, 32'h42b9c9fc, 32'hc1e92637};
test_label[878] = '{32'h4242be9d};
test_output[878] = '{32'h4230d55b};
/*############ DEBUG ############
test_input[7024:7031] = '{-71.8118423028, -52.07550248, -7.40311381342, 48.6861468901, 16.9531767753, 10.3252010467, 92.8945025765, -29.1436591813};
test_label[878] = '{48.6861468901};
test_output[878] = '{44.2083556864};
############ END DEBUG ############*/
test_input[7032:7039] = '{32'hc229e9fe, 32'h42460ac9, 32'hc28ac078, 32'hc293045f, 32'h41b96597, 32'hc2b273db, 32'h42366012, 32'hc0ef816c};
test_label[879] = '{32'h41b96597};
test_output[879] = '{32'h41d2d85a};
/*############ DEBUG ############
test_input[7032:7039] = '{-42.4785074996, 49.5105329191, -69.3759180354, -73.5085402867, 23.174603815, -89.2262766987, 45.5938188051, -7.48454859495};
test_label[879] = '{23.174603815};
test_output[879] = '{26.35563996};
############ END DEBUG ############*/
test_input[7040:7047] = '{32'hc276f3bf, 32'hc2114ead, 32'h411e1505, 32'h42c7b81d, 32'h42057e80, 32'h40ec7d96, 32'h4206b207, 32'h4160bbb1};
test_label[880] = '{32'hc276f3bf};
test_output[880] = '{32'h432198fe};
/*############ DEBUG ############
test_input[7040:7047] = '{-61.7380346718, -36.3268303745, 9.8801313545, 99.8595969035, 33.3735355772, 7.39033038821, 33.6738537446, 14.0458232008};
test_label[880] = '{-61.7380346718};
test_output[880] = '{161.597631575};
############ END DEBUG ############*/
test_input[7048:7055] = '{32'h4137a761, 32'h42c1da14, 32'hc253ef5f, 32'hc2958e40, 32'hc2c617eb, 32'hc1cdaf70, 32'hc257fa37, 32'hc2aa37ab};
test_label[881] = '{32'hc2958e40};
test_output[881] = '{32'h432bb42a};
/*############ DEBUG ############
test_input[7048:7055] = '{11.4783641584, 96.9259343341, -52.9837608898, -74.7778298266, -99.0467134683, -25.7106625111, -53.9943491045, -85.1087265409};
test_label[881] = '{-74.7778298266};
test_output[881] = '{171.703764161};
############ END DEBUG ############*/
test_input[7056:7063] = '{32'h4247df89, 32'hc2735d3f, 32'hc285fb10, 32'h4145957a, 32'h42c468cd, 32'hc1ed8e6d, 32'hc125236b, 32'h425f063c};
test_label[882] = '{32'hc1ed8e6d};
test_output[882] = '{32'h42ffcc68};
/*############ DEBUG ############
test_input[7056:7063] = '{49.9682952822, -60.8410624047, -66.9903569578, 12.3489928381, 98.2046895877, -29.6945433369, -10.3211465417, 55.7560886638};
test_label[882] = '{-29.6945433369};
test_output[882] = '{127.899232925};
############ END DEBUG ############*/
test_input[7064:7071] = '{32'hc276fcd6, 32'h4263a1bd, 32'hc1775935, 32'hc0cb44ef, 32'hc28baa3a, 32'h42573161, 32'hc290d56f, 32'hc2b44937};
test_label[883] = '{32'hc28baa3a};
test_output[883] = '{32'h42fd9171};
/*############ DEBUG ############
test_input[7064:7071] = '{-61.7469096507, 56.9079478503, -15.4592790074, -6.35216466156, -69.8324738256, 53.7982201498, -72.4168601, -90.1429963268};
test_label[883] = '{-69.8324738256};
test_output[883] = '{126.784068255};
############ END DEBUG ############*/
test_input[7072:7079] = '{32'h40bb78cd, 32'h4284b4b5, 32'h429b18d4, 32'h42c17980, 32'h4232da80, 32'hc1e043b0, 32'hc1a4fd47, 32'hbf73a797};
test_label[884] = '{32'hc1a4fd47};
test_output[884] = '{32'h42eab8d2};
/*############ DEBUG ############
test_input[7072:7079] = '{5.85849632476, 66.3529421706, 77.5484893053, 96.7373066647, 44.713380536, -28.0330497828, -20.6236702934, -0.951775961872};
test_label[884] = '{-20.6236702934};
test_output[884] = '{117.360976963};
############ END DEBUG ############*/
test_input[7080:7087] = '{32'h4210d8b1, 32'hc2402cd5, 32'h419564c4, 32'h4234f7fe, 32'h4268b579, 32'h42bc979f, 32'hc218dc68, 32'hc2c73844};
test_label[885] = '{32'h4268b579};
test_output[885] = '{32'h421079c6};
/*############ DEBUG ############
test_input[7080:7087] = '{36.211613884, -48.0437820425, 18.6742013569, 45.24218064, 58.1772195989, 94.2961380416, -38.2152417918, -99.6098912028};
test_label[885] = '{58.1772195989};
test_output[885] = '{36.1189184427};
############ END DEBUG ############*/
test_input[7088:7095] = '{32'h429b6d66, 32'h41f23d4f, 32'h42c4c9e6, 32'hc1de00ba, 32'hc0cfd478, 32'hc17f09cd, 32'h4174d2b6, 32'hc0b62fb1};
test_label[886] = '{32'h4174d2b6};
test_output[886] = '{32'h42a62f8f};
/*############ DEBUG ############
test_input[7088:7095] = '{77.713668574, 30.2799349324, 98.3943292345, -27.7503551654, -6.49468636492, -15.9398923414, 15.3014427095, -5.6933216233};
test_label[886] = '{15.3014427095};
test_output[886] = '{83.0928865261};
############ END DEBUG ############*/
test_input[7096:7103] = '{32'h42befc66, 32'hc29c2e20, 32'h3e9080df, 32'hc27a532b, 32'hc2bf27fd, 32'hc1a61882, 32'hc2b6c1e9, 32'h42a844d2};
test_label[887] = '{32'hc29c2e20};
test_output[887] = '{32'h432d9544};
/*############ DEBUG ############
test_input[7096:7103] = '{95.4929680547, -78.0900861567, 0.28223321357, -62.5812195378, -95.5781043097, -20.7619672163, -91.3787333175, 84.13441382};
test_label[887] = '{-78.0900861567};
test_output[887] = '{173.583065881};
############ END DEBUG ############*/
test_input[7104:7111] = '{32'hc1c9554d, 32'hc0cc1200, 32'h4244e6c8, 32'h41768036, 32'h427feceb, 32'hc16cc3f7, 32'hc158ab84, 32'h422cdd45};
test_label[888] = '{32'hc1c9554d};
test_output[888] = '{32'h42b24bc9};
/*############ DEBUG ############
test_input[7104:7111] = '{-25.1666508412, -6.37719720023, 49.2253738255, 15.4063010657, 63.9813636011, -14.7978426532, -13.541874382, 43.2160833033};
test_label[888] = '{-25.1666508412};
test_output[888] = '{89.1480148337};
############ END DEBUG ############*/
test_input[7112:7119] = '{32'hc266bf6e, 32'h41cc03ba, 32'hc0b791c5, 32'hc1306bf9, 32'h4298ecdf, 32'hc1a6750c, 32'hc1d8dcc8, 32'hc278a806};
test_label[889] = '{32'hc278a806};
test_output[889] = '{32'h430aa071};
/*############ DEBUG ############
test_input[7112:7119] = '{-57.6869440369, 25.5018191246, -5.73654435097, -11.0263605961, 76.4626385857, -20.8071514644, -27.1078026905, -62.1640860254};
test_label[889] = '{-62.1640860254};
test_output[889] = '{138.626724611};
############ END DEBUG ############*/
test_input[7120:7127] = '{32'h4185a070, 32'hc27284b6, 32'h42985b7b, 32'h422cf229, 32'hc1017270, 32'hc19c3c78, 32'hc25351c1, 32'h42c13ee7};
test_label[890] = '{32'h4185a070};
test_output[890] = '{32'h429fd6cb};
/*############ DEBUG ############
test_input[7120:7127] = '{16.7033381473, -60.6296022557, 76.1786749298, 43.2364827103, -8.09043925184, -19.5295265662, -52.8298372409, 96.6228525634};
test_label[890] = '{16.7033381473};
test_output[890] = '{79.9195144174};
############ END DEBUG ############*/
test_input[7128:7135] = '{32'hc088e18f, 32'hc1b4f385, 32'hc1fde099, 32'h424ae108, 32'h410e5543, 32'hc29dea99, 32'h428eac8a, 32'hc1fe4387};
test_label[891] = '{32'hc088e18f};
test_output[891] = '{32'h42973aa3};
/*############ DEBUG ############
test_input[7128:7135] = '{-4.27753378658, -22.6189060129, -31.7346662011, 50.7197552166, 8.89581601533, -78.9582022358, 71.336992913, -31.7829731604};
test_label[891] = '{-4.27753378658};
test_output[891] = '{75.6145267007};
############ END DEBUG ############*/
test_input[7136:7143] = '{32'h42abb3ab, 32'h42923dfe, 32'h41ed33f1, 32'hc211c535, 32'hc18e4b25, 32'hc2c19ad6, 32'h42450c09, 32'h42312d07};
test_label[892] = '{32'h42923dfe};
test_output[892] = '{32'h414bad6e};
/*############ DEBUG ############
test_input[7136:7143] = '{85.850916669, 73.1210785813, 29.6503620447, -36.4425841786, -17.7866919466, -96.8024136939, 49.2617533102, 44.2939710173};
test_label[892] = '{73.1210785813};
test_output[892] = '{12.7298410492};
############ END DEBUG ############*/
test_input[7144:7151] = '{32'h40c5032d, 32'hc27a3dab, 32'hc25cea11, 32'h42aaff98, 32'h4176fdb0, 32'h429d03e8, 32'hc2b992d1, 32'hc1d3f9b2};
test_label[893] = '{32'h429d03e8};
test_output[893] = '{32'h40dfc287};
/*############ DEBUG ############
test_input[7144:7151] = '{6.15663771787, -62.5602230399, -55.228578707, 85.4992034775, 15.4369356939, 78.5076267222, -92.7867516688, -26.4969208267};
test_label[893] = '{78.5076267222};
test_output[893] = '{6.99249592811};
############ END DEBUG ############*/
test_input[7152:7159] = '{32'hc19deddd, 32'h4198e31d, 32'h4231a195, 32'h41f4004a, 32'hc2a31142, 32'h421a97c7, 32'hc29d4fdb, 32'h41fc87b4};
test_label[894] = '{32'h4231a195};
test_output[894] = '{32'h3b4e81c4};
/*############ DEBUG ############
test_input[7152:7159] = '{-19.7411433958, 19.11089466, 44.4077932119, 30.5001411491, -81.5337078594, 38.6482193185, -78.6559679078, 31.5662610911};
test_label[894] = '{44.4077932119};
test_output[894] = '{0.00315104527896};
############ END DEBUG ############*/
test_input[7160:7167] = '{32'h428c2673, 32'hc14f6d27, 32'h428220dd, 32'h415a89df, 32'h428cad2b, 32'hc2597812, 32'h425e457e, 32'hc165a7a6};
test_label[895] = '{32'h428c2673};
test_output[895] = '{32'h3f561300};
/*############ DEBUG ############
test_input[7160:7167] = '{70.0750981288, -12.964148324, 65.0641894847, 13.6586596794, 70.3382155383, -54.3672576704, 55.5678645271, -14.3534301294};
test_label[895] = '{70.0750981288};
test_output[895] = '{0.836227438468};
############ END DEBUG ############*/
test_input[7168:7175] = '{32'h421b18ab, 32'h429682e8, 32'hc121b45a, 32'h421b38d4, 32'h4281a2e9, 32'hc2a37b34, 32'h42968385, 32'hc1c6ea82};
test_label[896] = '{32'hc2a37b34};
test_output[896] = '{32'h431db0a8};
/*############ DEBUG ############
test_input[7168:7175] = '{38.774089035, 75.2556743136, -10.1065312646, 38.8054979347, 64.8181829052, -81.7406303515, 75.2568741056, -24.8645049265};
test_label[896] = '{-81.7406303515};
test_output[896] = '{157.690066569};
############ END DEBUG ############*/
test_input[7176:7183] = '{32'h413adaae, 32'hc285efa3, 32'hc2ad63bd, 32'h41b8f269, 32'h427c9b6d, 32'h422ebff1, 32'hc29cdaa9, 32'h42781018};
test_label[897] = '{32'h42781018};
test_output[897] = '{32'h3fb50ecf};
/*############ DEBUG ############
test_input[7176:7183] = '{11.6783885134, -66.9680435125, -86.694797777, 23.1183645343, 63.1517831161, 43.6874410178, -78.4270695502, 62.0157183035};
test_label[897] = '{62.0157183035};
test_output[897] = '{1.41451443632};
############ END DEBUG ############*/
test_input[7184:7191] = '{32'hc2751023, 32'h426ff40a, 32'h41828804, 32'hc245feea, 32'h42b28b13, 32'hc29973f6, 32'h40b4911c, 32'hc2b39aed};
test_label[898] = '{32'h41828804};
test_output[898] = '{32'h4291e912};
/*############ DEBUG ############
test_input[7184:7191] = '{-61.2657603977, 59.9883177744, 16.3164147579, -49.4989404381, 89.2716328896, -76.7264844497, 5.64271377813, -89.8025926797};
test_label[898] = '{16.3164147579};
test_output[898] = '{72.9552181317};
############ END DEBUG ############*/
test_input[7192:7199] = '{32'hc25013ec, 32'hc1bd096d, 32'h42b6e8a4, 32'h42b89fae, 32'hc2adf075, 32'h42b1cc87, 32'hbebb5cd8, 32'h424f1797};
test_label[899] = '{32'h42b1cc87};
test_output[899] = '{32'h40727d7d};
/*############ DEBUG ############
test_input[7192:7199] = '{-52.0194558097, -23.6296021012, 91.4543752701, 92.3118707902, -86.9696428069, 88.8994682616, -0.365942708359, 51.773036945};
test_label[899] = '{88.8994682616};
test_output[899] = '{3.78890910658};
############ END DEBUG ############*/
test_input[7200:7207] = '{32'h42706892, 32'hc2ac99c6, 32'hc24ab158, 32'h42b65bba, 32'h42b26332, 32'hc243e795, 32'h40cc4f3a, 32'hc28e99a1};
test_label[900] = '{32'h42b65bba};
test_output[900] = '{32'h3e03c42c};
/*############ DEBUG ############
test_input[7200:7207] = '{60.1021202492, -86.3003368102, -50.6731879096, 91.1791510607, 89.1937380153, -48.9761559032, 6.38467134777, -71.3000592925};
test_label[900] = '{91.1791510607};
test_output[900] = '{0.128678030328};
############ END DEBUG ############*/
test_input[7208:7215] = '{32'h4246e7e8, 32'hc0db75cc, 32'h41263d35, 32'hc2ba9826, 32'hc2c0b38d, 32'h42b7c4a6, 32'h427797c6, 32'hc258dd0d};
test_label[901] = '{32'hc2ba9826};
test_output[901] = '{32'h43392e66};
/*############ DEBUG ############
test_input[7208:7215] = '{49.726469858, -6.85812966567, 10.3899430321, -93.2971661459, -96.3506881205, 91.884079505, 61.8982179489, -54.2158706936};
test_label[901] = '{-93.2971661459};
test_output[901] = '{185.181245651};
############ END DEBUG ############*/
test_input[7216:7223] = '{32'h4191334e, 32'hc258374f, 32'hc1f19e3b, 32'hc26df479, 32'h42a76095, 32'hc27becd6, 32'hc28ae441, 32'hc2950fb7};
test_label[902] = '{32'h42a76095};
test_output[902] = '{32'h80000000};
/*############ DEBUG ############
test_input[7216:7223] = '{18.1500510886, -54.0540111621, -30.2022615913, -59.4887421344, 83.6886370339, -62.9812850659, -69.4458105954, -74.5306921138};
test_label[902] = '{83.6886370339};
test_output[902] = '{-0.0};
############ END DEBUG ############*/
test_input[7224:7231] = '{32'h4299d0b9, 32'h41bcdb20, 32'h42aed8a3, 32'hc23b7457, 32'h3ee0e7cc, 32'h41d431e1, 32'h42b45d2e, 32'h42afbba2};
test_label[903] = '{32'h3ee0e7cc};
test_output[903] = '{32'h42b3c92e};
/*############ DEBUG ############
test_input[7224:7231] = '{76.907664602, 23.6069953915, 87.4231181324, -46.8636116782, 0.439268465052, 26.5243558746, 90.1819883388, 87.8664740689};
test_label[903] = '{0.439268465052};
test_output[903] = '{89.8929317535};
############ END DEBUG ############*/
test_input[7232:7239] = '{32'hc184b1da, 32'h42ac5ce3, 32'h41f4fb43, 32'h424dd827, 32'h4208b2c1, 32'hc2741282, 32'hc2be3666, 32'hc232074d};
test_label[904] = '{32'h424dd827};
test_output[904] = '{32'h420ae19f};
/*############ DEBUG ############
test_input[7232:7239] = '{-16.5868415698, 86.181417477, 30.6226857547, 51.4610845967, 34.1745636431, -61.0180738953, -95.1062443233, -44.507128416};
test_label[904] = '{51.4610845967};
test_output[904] = '{34.7203328803};
############ END DEBUG ############*/
test_input[7240:7247] = '{32'hc1d6f428, 32'hc25dbda7, 32'hc28f4dee, 32'hc2838af7, 32'hc2b7dc14, 32'h42763792, 32'hc29325a7, 32'hc2c0ce28};
test_label[905] = '{32'hc28f4dee};
test_output[905] = '{32'h430534db};
/*############ DEBUG ############
test_input[7240:7247] = '{-26.8692173835, -55.43520851, -71.6522053092, -65.7714186441, -91.9298434655, 61.5542668024, -73.5735372932, -96.402646771};
test_label[905] = '{-71.6522053092};
test_output[905] = '{133.206472112};
############ END DEBUG ############*/
test_input[7248:7255] = '{32'hc1ff15ea, 32'h420bb2ac, 32'h420fc0d6, 32'hc2c77651, 32'h4261bedd, 32'hc1ca057f, 32'h4192451b, 32'hc1f6e17b};
test_label[906] = '{32'h4192451b};
test_output[906] = '{32'h42189c50};
/*############ DEBUG ############
test_input[7248:7255] = '{-31.8857001138, 34.9244853953, 35.9383177002, -99.7310868326, 56.4363904051, -25.2526828984, 18.2837422829, -30.8600972329};
test_label[906] = '{18.2837422829};
test_output[906] = '{38.1526481239};
############ END DEBUG ############*/
test_input[7256:7263] = '{32'h424ddca2, 32'h41cbf19e, 32'h420ad76f, 32'h3fd526b8, 32'hc2b1eef8, 32'hc22ba1bf, 32'h429dcb87, 32'h42535a33};
test_label[907] = '{32'h42535a33};
test_output[907] = '{32'h41d079b6};
/*############ DEBUG ############
test_input[7256:7263] = '{51.4654621675, 25.4929771241, 34.7103850224, 1.66524415481, -88.9667360314, -42.9079532834, 78.8975129729, 52.8380843154};
test_label[907] = '{52.8380843154};
test_output[907] = '{26.0594286574};
############ END DEBUG ############*/
test_input[7264:7271] = '{32'hc298023d, 32'h42a4d181, 32'h424111d1, 32'h407c55fa, 32'h4282eecd, 32'h4154fd01, 32'hbe994f15, 32'hc284afcd};
test_label[908] = '{32'hc284afcd};
test_output[908] = '{32'h4314c0a7};
/*############ DEBUG ############
test_input[7264:7271] = '{-76.0043711764, 82.4091855185, 48.2674005421, 3.94274759124, 65.4664105408, 13.3117683141, -0.299431484246, -66.3433640934};
test_label[908] = '{-66.3433640934};
test_output[908] = '{148.752549656};
############ END DEBUG ############*/
test_input[7272:7279] = '{32'hc295e8e0, 32'hc29cf2e3, 32'hc24bd8a1, 32'hc17ec886, 32'hc2114363, 32'hc1b8917b, 32'h422ba10b, 32'h4182f08b};
test_label[909] = '{32'h4182f08b};
test_output[909] = '{32'h41d4518a};
/*############ DEBUG ############
test_input[7272:7279] = '{-74.954831058, -78.4743912423, -50.9615512972, -15.9239560544, -36.3158089971, -23.0710348356, 42.9072668861, 16.3674527936};
test_label[909] = '{16.3674527936};
test_output[909] = '{26.5398140925};
############ END DEBUG ############*/
test_input[7280:7287] = '{32'h4232ee7b, 32'h426818ca, 32'h421dcdfd, 32'h41256ce7, 32'h42b7d162, 32'h42c04f15, 32'h428dbcac, 32'h42c10a95};
test_label[910] = '{32'h42c10a95};
test_output[910] = '{32'h3f085608};
/*############ DEBUG ############
test_input[7280:7287] = '{44.7328912997, 58.0242073164, 39.4511599658, 10.3390876847, 91.9089518163, 96.1544595764, 70.8684971887, 96.5206697265};
test_label[910] = '{96.5206697265};
test_output[910] = '{0.532562739594};
############ END DEBUG ############*/
test_input[7288:7295] = '{32'h3f4e5938, 32'h40e4e698, 32'hc29f38af, 32'hc2b06cdf, 32'hc28104c9, 32'hc1c846c1, 32'h41061111, 32'h40e687cd};
test_label[911] = '{32'h41061111};
test_output[911] = '{32'h3ef18696};
/*############ DEBUG ############
test_input[7288:7295] = '{0.806048860849, 7.15314879553, -79.6107129207, -88.2126411466, -64.509344242, -25.0345486424, 8.37916635406, 7.20407714648};
test_label[911] = '{8.37916635406};
test_output[911] = '{0.471729923284};
############ END DEBUG ############*/
test_input[7296:7303] = '{32'h40626ddc, 32'h42a99b3f, 32'h413f7316, 32'h4243169a, 32'hc1c17b2c, 32'hc2a4b759, 32'h42ad40e5, 32'h41d1c600};
test_label[912] = '{32'h42ad40e5};
test_output[912] = '{32'h3e1943ba};
/*############ DEBUG ############
test_input[7296:7303] = '{3.53795517817, 84.8032127247, 11.9655967994, 48.7720727742, -24.1851431217, -82.3580990505, 86.6267495087, 26.221679965};
test_label[912] = '{86.6267495087};
test_output[912] = '{0.149672421409};
############ END DEBUG ############*/
test_input[7304:7311] = '{32'h41eb46ea, 32'h4164da39, 32'hc145c05f, 32'h42198735, 32'hc2b34937, 32'h42bcbcd6, 32'hc2374970, 32'hc291db18};
test_label[913] = '{32'h4164da39};
test_output[913] = '{32'h42a0218e};
/*############ DEBUG ############
test_input[7304:7311] = '{29.4096263178, 14.303277305, -12.3594654117, 38.3820390392, -89.6430004106, 94.368817157, -45.8217176008, -72.9279198835};
test_label[913] = '{14.303277305};
test_output[913] = '{80.065539852};
############ END DEBUG ############*/
test_input[7312:7319] = '{32'h4137bf29, 32'h4255eb02, 32'h414c6d3a, 32'h40656c49, 32'hc1e0702a, 32'h4238ddeb, 32'h42a4d441, 32'hc2088397};
test_label[914] = '{32'h4137bf29};
test_output[914] = '{32'h428ddc5c};
/*############ DEBUG ############
test_input[7312:7319] = '{11.4841702697, 53.4795009395, 12.7766671177, 3.58473430387, -28.0547678249, 46.2167169697, 82.4145609826, -34.128504214};
test_label[914] = '{11.4841702697};
test_output[914] = '{70.9303907128};
############ END DEBUG ############*/
test_input[7320:7327] = '{32'h41d580a1, 32'h4218ec2a, 32'h40d13ae6, 32'h3ec723f0, 32'hc294adc5, 32'hc1ed5dd2, 32'h423193ec, 32'hc2a7e84a};
test_label[915] = '{32'hc2a7e84a};
test_output[915] = '{32'h430059aa};
/*############ DEBUG ############
test_input[7320:7327] = '{26.6878076482, 38.23062804, 6.53843973658, 0.388946044358, -74.3393911874, -29.670810128, 44.3944552623, -83.9536869367};
test_label[915] = '{-83.9536869367};
test_output[915] = '{128.350244193};
############ END DEBUG ############*/
test_input[7328:7335] = '{32'h41ca6b8c, 32'h423d7b9c, 32'hc0e5db87, 32'h41771cec, 32'h42197f50, 32'h400ea7ec, 32'h41fc7b92, 32'hc1ec9766};
test_label[916] = '{32'h42197f50};
test_output[916] = '{32'h410ff1b0};
/*############ DEBUG ############
test_input[7328:7335] = '{25.3025136037, 47.3707106547, -7.18304766891, 15.4445608315, 38.3743286392, 2.22899914066, 31.560336843, -29.573925344};
test_label[916] = '{38.3743286392};
test_output[916] = '{8.99650600115};
############ END DEBUG ############*/
test_input[7336:7343] = '{32'h42115288, 32'h415d374b, 32'hc108a664, 32'h42074b42, 32'hc2a58417, 32'hc1b8463e, 32'h4295bc62, 32'h42a9894c};
test_label[917] = '{32'h415d374b};
test_output[917] = '{32'h428de269};
/*############ DEBUG ############
test_input[7336:7343] = '{36.3305979281, 13.8259990141, -8.54062288586, 33.8234922428, -82.7579861479, -23.0342982261, 74.8679357754, 84.7681583555};
test_label[917] = '{13.8259990141};
test_output[917] = '{70.9422095037};
############ END DEBUG ############*/
test_input[7344:7351] = '{32'hc2b1b7cf, 32'hc2898568, 32'hc21c6e52, 32'hc2598228, 32'hc2565a91, 32'hc0524660, 32'hc208046c, 32'h42a09e60};
test_label[918] = '{32'hc2b1b7cf};
test_output[918] = '{32'h43292b18};
/*############ DEBUG ############
test_input[7344:7351] = '{-88.8590040533, -68.7605597165, -39.107734761, -54.3771044019, -53.5884428284, -3.28554543199, -34.0043197146, 80.3093284547};
test_label[918] = '{-88.8590040533};
test_output[918] = '{169.168332508};
############ END DEBUG ############*/
test_input[7352:7359] = '{32'h425c5f50, 32'h4130820f, 32'hc03770c2, 32'h41b5ab2f, 32'h4282f21d, 32'hc2c2f4f4, 32'hc243a51c, 32'hc2a4b686};
test_label[919] = '{32'h4130820f};
test_output[919] = '{32'h4259c3bf};
/*############ DEBUG ############
test_input[7352:7359] = '{55.0930790291, 11.0317524277, -2.86625723475, 22.7085850515, 65.4728784893, -97.4784227236, -48.9112395822, -82.3564927418};
test_label[919] = '{11.0317524277};
test_output[919] = '{54.4411571147};
############ END DEBUG ############*/
test_input[7360:7367] = '{32'h42170349, 32'h4232de44, 32'h412ea6f9, 32'hc205c1e5, 32'hc26aeef6, 32'hc27c1878, 32'hc16367f6, 32'hc18b1252};
test_label[920] = '{32'hc18b1252};
test_output[920] = '{32'h42786864};
/*############ DEBUG ############
test_input[7360:7367] = '{37.7532090032, 44.7170559806, 10.9157649654, -33.43935184, -58.7333584307, -63.0238965882, -14.212880687, -17.3839447051};
test_label[920] = '{-17.3839447051};
test_output[920] = '{62.1019456914};
############ END DEBUG ############*/
test_input[7368:7375] = '{32'hc2695800, 32'hbf359b07, 32'h426802a3, 32'h42919ced, 32'h4206153b, 32'h428a89ab, 32'h42831c5f, 32'h423a43a9};
test_label[921] = '{32'h4206153b};
test_output[921] = '{32'h421d42af};
/*############ DEBUG ############
test_input[7368:7375] = '{-58.3359369028, -0.70939677215, 58.0025737921, 72.8064945803, 33.5207310577, 69.2688814546, 65.5554142144, 46.566072496};
test_label[921] = '{33.5207310577};
test_output[921] = '{39.3151207906};
############ END DEBUG ############*/
test_input[7376:7383] = '{32'hc2b5651b, 32'h419f3ae2, 32'hc2c72d8a, 32'h42846c54, 32'hc264f228, 32'hc2967d52, 32'hc2486282, 32'hc237e199};
test_label[922] = '{32'hc237e199};
test_output[922] = '{32'h42e05d20};
/*############ DEBUG ############
test_input[7376:7383] = '{-90.6974694965, 19.9037508714, -99.5889403959, 66.2115766237, -57.2364809555, -75.2447638697, -50.096198783, -45.9703100043};
test_label[922] = '{-45.9703100043};
test_output[922] = '{112.181886628};
############ END DEBUG ############*/
test_input[7384:7391] = '{32'hc2bd696f, 32'hc26c36ab, 32'h42c121f6, 32'h423a051c, 32'hc1bf29ce, 32'h421d4f46, 32'h4259df79, 32'hc2c10ef7};
test_label[923] = '{32'h4259df79};
test_output[923] = '{32'h42286473};
/*############ DEBUG ############
test_input[7384:7391] = '{-94.7059249481, -59.0533883162, 96.56633133, 46.5049888772, -23.8954121709, 39.3274154572, 54.4682363323, -96.5292275905};
test_label[923] = '{54.4682363323};
test_output[923] = '{42.0980949977};
############ END DEBUG ############*/
test_input[7392:7399] = '{32'hc24a9bf5, 32'h424dcba3, 32'hc2c483e7, 32'hc18857b3, 32'hc2a0c7cf, 32'h4104eabe, 32'h4287d721, 32'h41ddbf70};
test_label[924] = '{32'hc2c483e7};
test_output[924] = '{32'h43262d84};
/*############ DEBUG ############
test_input[7392:7399] = '{-50.6523008568, 51.4488621809, -98.2576227416, -17.0428210405, -80.3902487935, 8.30731018383, 67.9201757605, 27.7184757841};
test_label[924] = '{-98.2576227416};
test_output[924] = '{166.177798572};
############ END DEBUG ############*/
test_input[7400:7407] = '{32'hbfabf247, 32'hc260c97c, 32'hc20b00d7, 32'h41b289a2, 32'hc21096f1, 32'h42a13206, 32'h41f56408, 32'hc16f89c1};
test_label[925] = '{32'hc21096f1};
test_output[925] = '{32'h42e97d7e};
/*############ DEBUG ############
test_input[7400:7407] = '{-1.34333121131, -56.1967622577, -34.7508208551, 22.3172027752, -36.1474034865, 80.5977016533, 30.673843554, -14.9711310556};
test_label[925] = '{-36.1474034865};
test_output[925] = '{116.74510514};
############ END DEBUG ############*/
test_input[7408:7415] = '{32'hc2ac8d79, 32'hc2adbf70, 32'h427cfb82, 32'hc217103a, 32'h42b3ca93, 32'hc1753eb3, 32'hc28be65a, 32'hc2580ece};
test_label[926] = '{32'hc2580ece};
test_output[926] = '{32'h430fe8fd};
/*############ DEBUG ############
test_input[7408:7415] = '{-86.2763157359, -86.8738982896, 63.2456146918, -37.7658462475, 89.8956541941, -15.3278072196, -69.9499084222, -54.0144589564};
test_label[926] = '{-54.0144589564};
test_output[926] = '{143.91011315};
############ END DEBUG ############*/
test_input[7416:7423] = '{32'h422f9257, 32'h42b5c4bf, 32'h410ab297, 32'h418ae3d5, 32'hc02debdf, 32'h4230173e, 32'hc243df71, 32'h428e0be3};
test_label[927] = '{32'h422f9257};
test_output[927] = '{32'h423bf726};
/*############ DEBUG ############
test_input[7416:7423] = '{43.8929110507, 90.8842661061, 8.66860116606, 17.3612465071, -2.71752133811, 44.0226969851, -48.9682033588, 71.0232132964};
test_label[927] = '{43.8929110507};
test_output[927] = '{46.9913550578};
############ END DEBUG ############*/
test_input[7424:7431] = '{32'h42c67a71, 32'h4198d9d8, 32'hc20a01e7, 32'h4286b5d1, 32'h425ca5bb, 32'h423c81ec, 32'h4088a76a, 32'hc29778ea};
test_label[928] = '{32'h423c81ec};
test_output[928] = '{32'h425072f6};
/*############ DEBUG ############
test_input[7424:7431] = '{99.2391425227, 19.1063684621, -34.5018596607, 67.3551068793, 55.1618459213, 47.1268768675, 4.27043616006, -75.736157282};
test_label[928] = '{47.1268768675};
test_output[928] = '{52.1122656553};
############ END DEBUG ############*/
test_input[7432:7439] = '{32'hc080aac8, 32'hc18cea17, 32'h42300989, 32'h429692e8, 32'hc2856922, 32'hc2ab459b, 32'hc282a6d8, 32'hc24be1e8};
test_label[929] = '{32'hc2856922};
test_output[929] = '{32'h430dfe05};
/*############ DEBUG ############
test_input[7432:7439] = '{-4.02084723349, -17.6143016309, 44.0093113908, 75.2869239417, -66.7053372781, -85.6359497321, -65.3258633309, -50.9706127007};
test_label[929] = '{-66.7053372781};
test_output[929] = '{141.99226122};
############ END DEBUG ############*/
test_input[7440:7447] = '{32'h423d458f, 32'hc2875465, 32'h41da8d1f, 32'h42b2755d, 32'hc21b36c7, 32'h4259a28c, 32'h420ae395, 32'hc2c35a0a};
test_label[930] = '{32'hc2c35a0a};
test_output[930] = '{32'h433ae7b3};
/*############ DEBUG ############
test_input[7440:7447] = '{47.3179274482, -67.6648329522, 27.3189062606, 89.2292246876, -38.8034943113, 54.408738283, 34.7222470778, -97.675854468};
test_label[930] = '{-97.675854468};
test_output[930] = '{186.905079156};
############ END DEBUG ############*/
test_input[7448:7455] = '{32'hc0bc6b44, 32'h429e2538, 32'h42ab5a16, 32'hc15c5f29, 32'h428fd492, 32'h4206bc6d, 32'hbf60fce6, 32'h42be1499};
test_label[931] = '{32'hc15c5f29};
test_output[931] = '{32'h42d9a089};
/*############ DEBUG ############
test_input[7448:7455] = '{-5.88809384092, 79.0726893338, 85.6759479559, -13.7732326149, 71.9151733689, 33.6840082233, -0.878858953111, 95.0402288376};
test_label[931] = '{-13.7732326149};
test_output[931] = '{108.813547297};
############ END DEBUG ############*/
test_input[7456:7463] = '{32'hc2bb0028, 32'h41a3ac2f, 32'h425d72f1, 32'hc2bfdaba, 32'hc24920ec, 32'hc238d3a9, 32'h42ba3623, 32'h4223bca7};
test_label[932] = '{32'hc2bfdaba};
test_output[932] = '{32'h433d086e};
/*############ DEBUG ############
test_input[7456:7463] = '{-93.500306179, 20.4590733963, 55.3622480385, -95.9271994325, -50.2821484235, -46.206699854, 93.1057348924, 40.9342309163};
test_label[932] = '{-95.9271994325};
test_output[932] = '{189.032934325};
############ END DEBUG ############*/
test_input[7464:7471] = '{32'h42b88084, 32'h42af4d68, 32'hc2bc43a6, 32'h41ffbddf, 32'hc2052508, 32'hc2c5fd73, 32'hc1fe6735, 32'hc1d33c8f};
test_label[933] = '{32'h41ffbddf};
test_output[933] = '{32'h42712c58};
/*############ DEBUG ############
test_input[7464:7471] = '{92.2510093198, 87.6511838095, -94.1321253892, 31.9677096162, -33.2861631172, -98.9950212169, -31.8003934037, -26.4045702376};
test_label[933] = '{31.9677096162};
test_output[933] = '{60.2933030923};
############ END DEBUG ############*/
test_input[7472:7479] = '{32'h41cb8b2b, 32'h3f7bf656, 32'hc2694951, 32'hc2b33144, 32'h4291370d, 32'hc1cca24b, 32'h428150bd, 32'h42c43637};
test_label[934] = '{32'hc2694951};
test_output[934] = '{32'h431c6d6f};
/*############ DEBUG ############
test_input[7472:7479] = '{25.4429529033, 0.984227550154, -58.3215970618, -89.5962207273, 72.6075197878, -25.5792451765, 64.6576930459, 98.1058853152};
test_label[934] = '{-58.3215970618};
test_output[934] = '{156.427482377};
############ END DEBUG ############*/
test_input[7480:7487] = '{32'hc1c076cc, 32'h429dac1f, 32'h429e6eb8, 32'h41e01310, 32'h4231aee1, 32'hc2beb79b, 32'hc251265c, 32'hc0a45fe0};
test_label[935] = '{32'h429dac1f};
test_output[935] = '{32'h3f66b0d6};
/*############ DEBUG ############
test_input[7480:7487] = '{-24.0580063148, 78.8361722478, 79.2162500149, 28.009306985, 44.4207810742, -95.3586066331, -52.2874618436, -5.1367036594};
test_label[935] = '{78.8361722478};
test_output[935] = '{0.90113579836};
############ END DEBUG ############*/
test_input[7488:7495] = '{32'h4114f5e6, 32'hc234821e, 32'h424f7b2d, 32'hc28899e4, 32'h429b33f7, 32'hc2af0071, 32'hc126f2f3, 32'hc28deb45};
test_label[936] = '{32'h429b33f7};
test_output[936] = '{32'h2ceb3200};
/*############ DEBUG ############
test_input[7488:7495] = '{9.31003415472, -45.1270668698, 51.8702871641, -68.3005657028, 77.6014922129, -87.5008600707, -10.4343136759, -70.9595113945};
test_label[936] = '{77.6014922129};
test_output[936] = '{6.68465283129e-12};
############ END DEBUG ############*/
test_input[7496:7503] = '{32'hc1f23f70, 32'hc1b332c3, 32'h425128a0, 32'h41e0b3e2, 32'h41d72a88, 32'h42661406, 32'hc2b61519, 32'h421e79d3};
test_label[937] = '{32'hc2b61519};
test_output[937] = '{32'h431490ec};
/*############ DEBUG ############
test_input[7496:7503] = '{-30.2809758144, -22.3997851657, 52.2896742417, 28.0878326322, 26.8957668032, 57.5195543289, -91.0412059841, 39.6189693386};
test_label[937] = '{-91.0412059841};
test_output[937] = '{148.566100214};
############ END DEBUG ############*/
test_input[7504:7511] = '{32'h42adef6f, 32'h42941a3a, 32'hc26e6a57, 32'hc1ce7703, 32'h420a823c, 32'hc0d3ee3b, 32'hc1b34538, 32'hc269bf02};
test_label[938] = '{32'h42941a3a};
test_output[938] = '{32'h414ea9a8};
/*############ DEBUG ############
test_input[7504:7511] = '{86.967641131, 74.0512236266, -59.6038482627, -25.8081104723, 34.627180962, -6.62283102919, -22.4087991224, -58.4365316718};
test_label[938] = '{74.0512236266};
test_output[938] = '{12.9164199618};
############ END DEBUG ############*/
test_input[7512:7519] = '{32'h42b09c84, 32'hc2a138ad, 32'h412edc09, 32'h423c7941, 32'hc29fd3d3, 32'hc29ef6f2, 32'hc2af34c8, 32'hc2ad6ac1};
test_label[939] = '{32'h423c7941};
test_output[939] = '{32'h4224bfc7};
/*############ DEBUG ############
test_input[7512:7519] = '{88.3056933108, -80.6106976602, 10.9287199087, 47.118411077, -79.9137191979, -79.4823175208, -87.603091961, -86.7085054722};
test_label[939] = '{47.118411077};
test_output[939] = '{41.1872822338};
############ END DEBUG ############*/
test_input[7520:7527] = '{32'hc2aece6f, 32'hc161d28c, 32'h422a5577, 32'hc2c5a7a9, 32'hc2887df9, 32'hc1f3bfc9, 32'hc242af84, 32'hc0a14e77};
test_label[940] = '{32'hc242af84};
test_output[940] = '{32'h42b6827e};
/*############ DEBUG ############
test_input[7520:7527] = '{-87.4031894366, -14.1139034284, 42.5834630518, -98.8274592936, -68.2460378335, -30.4686449075, -48.6714026046, -5.0408282396};
test_label[940] = '{-48.6714026046};
test_output[940] = '{91.2548656564};
############ END DEBUG ############*/
test_input[7528:7535] = '{32'h418dc97b, 32'h41fec3b7, 32'hc07ca4d6, 32'hc298a08f, 32'h4279ab0f, 32'hc262342f, 32'hc2920a75, 32'hc1ae8f90};
test_label[941] = '{32'hc262342f};
test_output[941] = '{32'h42edef9f};
/*############ DEBUG ############
test_input[7528:7535] = '{17.7233800526, 31.8455633343, -3.94756087836, -76.31359048, 62.4170503584, -56.5509619492, -73.0204259057, -21.8200986745};
test_label[941] = '{-56.5509619492};
test_output[941] = '{118.968012308};
############ END DEBUG ############*/
test_input[7536:7543] = '{32'hc1c808b4, 32'hc2aae903, 32'hc0099069, 32'h41f3b8d4, 32'hc1f7462e, 32'h42c2af1d, 32'h417b7533, 32'h4273324a};
test_label[942] = '{32'h417b7533};
test_output[942] = '{32'h42a34076};
/*############ DEBUG ############
test_input[7536:7543] = '{-25.0042498301, -85.4551048141, -2.14943920111, 30.4652478354, -30.9092680622, 97.3420169292, 15.716113338, 60.7991099571};
test_label[942] = '{15.716113338};
test_output[942] = '{81.6259035912};
############ END DEBUG ############*/
test_input[7544:7551] = '{32'hc29f26c9, 32'hc297da10, 32'h41ce5a38, 32'hc2b95e22, 32'hc1918199, 32'h42bbaf07, 32'h413ada97, 32'h406a22e0};
test_label[943] = '{32'hc29f26c9};
test_output[943] = '{32'h432d6ae8};
/*############ DEBUG ############
test_input[7544:7551] = '{-79.5757517993, -75.9259038002, 25.7940513374, -92.6838541394, -18.1882803777, 93.8418509108, 11.6783662665, 3.65837858244};
test_label[943] = '{-79.5757517993};
test_output[943] = '{173.41760271};
############ END DEBUG ############*/
test_input[7552:7559] = '{32'h429bdc0b, 32'h427a2449, 32'hc1a0c02e, 32'hc1d427c2, 32'hc2b0855e, 32'h41e11d86, 32'hc2a79f4f, 32'h40f407e7};
test_label[944] = '{32'h429bdc0b};
test_output[944] = '{32'h345d6c5d};
/*############ DEBUG ############
test_input[7552:7559] = '{77.9297744188, 62.5354353543, -20.0938367917, -26.5194128732, -88.2604811247, 28.1394159347, -83.8111464531, 7.62596463031};
test_label[944] = '{77.9297744188};
test_output[944] = '{2.06216516809e-07};
############ END DEBUG ############*/
test_input[7560:7567] = '{32'hc2ba5cbe, 32'h42be7d4a, 32'hc1c5248c, 32'hc2147064, 32'hc2bfe3ae, 32'hc1b2872f, 32'hc204eb70, 32'hc28b57e4};
test_label[945] = '{32'hc2147064};
test_output[945] = '{32'h43045abe};
/*############ DEBUG ############
test_input[7560:7567] = '{-93.1811334949, 95.24470624, -24.6428442425, -37.1097558179, -95.9446881322, -22.3160067882, -33.2299210277, -69.6716615843};
test_label[945] = '{-37.1097558179};
test_output[945] = '{132.354462058};
############ END DEBUG ############*/
test_input[7568:7575] = '{32'hc05afa0b, 32'h422f2f7a, 32'h42c0eb59, 32'h4296a6b5, 32'h423e3679, 32'h429afaf9, 32'h416ab28e, 32'h429e3a7a};
test_label[946] = '{32'h422f2f7a};
test_output[946] = '{32'h4252a738};
/*############ DEBUG ############
test_input[7568:7575] = '{-3.42151132228, 43.7963628404, 96.4596624289, 75.325596137, 47.5531952826, 77.4901776124, 14.6685923432, 79.1142151359};
test_label[946] = '{43.7963628404};
test_output[946] = '{52.6632996242};
############ END DEBUG ############*/
test_input[7576:7583] = '{32'hc185aed0, 32'h428c6b1f, 32'hc2c5a90e, 32'hc282449a, 32'hc28d8cc0, 32'h42167cd4, 32'hc27a0cc4, 32'h42c105e6};
test_label[947] = '{32'hc27a0cc4};
test_output[947] = '{32'h431f0624};
/*############ DEBUG ############
test_input[7576:7583] = '{-16.7103573148, 70.2092245013, -98.8301814425, -65.1339858927, -70.7748997418, 37.6219026512, -62.5124667231, 96.5115175144};
test_label[947] = '{-62.5124667231};
test_output[947] = '{159.023984238};
############ END DEBUG ############*/
test_input[7584:7591] = '{32'h42a2f619, 32'h41d9affb, 32'h427dadf6, 32'hc291bef8, 32'hc214a199, 32'h4160d3c3, 32'h429e5965, 32'hc19b7cdb};
test_label[948] = '{32'h41d9affb};
test_output[948] = '{32'h4259757b};
/*############ DEBUG ############
test_input[7584:7591] = '{81.4806606425, 27.2109278918, 63.419885519, -72.8729876635, -37.1578114195, 14.0516994236, 79.1745952263, -19.4359650168};
test_label[948] = '{27.2109278918};
test_output[948] = '{54.3647270506};
############ END DEBUG ############*/
test_input[7592:7599] = '{32'hc1c87dbf, 32'hc2b41919, 32'hc19a5c02, 32'h42b8f2a8, 32'h425af607, 32'h425c1e17, 32'hc2a917e4, 32'h42954fb9};
test_label[949] = '{32'h42954fb9};
test_output[949] = '{32'h418e8bbd};
/*############ DEBUG ############
test_input[7592:7599] = '{-25.0614001953, -90.0490161126, -19.2949253061, 92.4739394979, 54.7402628695, 55.0293842569, -84.5466619513, 74.6557079139};
test_label[949] = '{74.6557079139};
test_output[949] = '{17.8182316023};
############ END DEBUG ############*/
test_input[7600:7607] = '{32'h4284f6db, 32'h42b8fa2c, 32'h4223708d, 32'hc25e401e, 32'hc27a275d, 32'h42b33b6e, 32'h42153e39, 32'h41e1b120};
test_label[950] = '{32'h4284f6db};
test_output[950] = '{32'h41d07dec};
/*############ DEBUG ############
test_input[7600:7607] = '{66.4821433179, 92.4886151952, 40.8599128153, -55.5626126284, -62.5384403875, 89.6160735371, 37.3107648936, 28.2114869332};
test_label[950] = '{66.4821433179};
test_output[950] = '{26.061485493};
############ END DEBUG ############*/
test_input[7608:7615] = '{32'h42b74ae5, 32'h42908f3f, 32'h409cf4c6, 32'hc259b752, 32'h41b02a36, 32'h425f4126, 32'h42c51b87, 32'h40af34c6};
test_label[951] = '{32'h409cf4c6};
test_output[951] = '{32'h42bb4cbe};
/*############ DEBUG ############
test_input[7608:7615] = '{91.6462751634, 72.2797753112, 4.90487941542, -54.4290244079, 22.0206099451, 55.8136221327, 98.5537653112, 5.47519197004};
test_label[951] = '{4.90487941542};
test_output[951] = '{93.6498856611};
############ END DEBUG ############*/
test_input[7616:7623] = '{32'h42692b78, 32'h42916b66, 32'hc261eb89, 32'h41f13a48, 32'hbfac3a1f, 32'h41e77008, 32'h40fbc7fe, 32'hc1b9066f};
test_label[952] = '{32'h42692b78};
test_output[952] = '{32'h4166ad51};
/*############ DEBUG ############
test_input[7616:7623] = '{58.2924492478, 72.7097619429, -56.4800150516, 30.1534580263, -1.34552369419, 28.9297034214, 7.86816313103, -23.1281420483};
test_label[952] = '{58.2924492478};
test_output[952] = '{14.417313243};
############ END DEBUG ############*/
test_input[7624:7631] = '{32'hc2b4b82d, 32'h42bf7bef, 32'hc283a59f, 32'hc261461a, 32'h42278d30, 32'h41901bf4, 32'h426743bb, 32'h42b31510};
test_label[953] = '{32'h42b31510};
test_output[953] = '{32'h40c67e8f};
/*############ DEBUG ############
test_input[7624:7631] = '{-90.3597148791, 95.742058895, -65.8234807328, -56.3184575488, 41.8878765657, 18.0136485365, 57.8161412014, 89.5411354681};
test_label[953] = '{89.5411354681};
test_output[953] = '{6.20294893166};
############ END DEBUG ############*/
test_input[7632:7639] = '{32'h42515190, 32'hc155b067, 32'hc211ecea, 32'hc1f43cad, 32'h4224d8c2, 32'h4180b426, 32'h40ff8172, 32'h41ed8a82};
test_label[954] = '{32'hc1f43cad};
test_output[954] = '{32'h42a5b7f5};
/*############ DEBUG ############
test_input[7632:7639] = '{52.3296500957, -13.3555670892, -36.4813600088, -30.5296263738, 41.2116793789, 16.0879628369, 7.9845511924, 29.6926316726};
test_label[954] = '{-30.5296263738};
test_output[954] = '{82.8592913127};
############ END DEBUG ############*/
test_input[7640:7647] = '{32'hc21914d0, 32'h4252d4d3, 32'h42391fdd, 32'hc25400b8, 32'hc06057c9, 32'hc290e3e8, 32'hc185bbd3, 32'h40bc3adf};
test_label[955] = '{32'hc21914d0};
test_output[955] = '{32'h42b5f5a6};
/*############ DEBUG ############
test_input[7640:7647] = '{-38.2703247767, 52.707837187, 46.2811173984, -53.0007011528, -3.50535808652, -72.4451291528, -16.7167105949, 5.88218618798};
test_label[955] = '{-38.2703247767};
test_output[955] = '{90.9797784052};
############ END DEBUG ############*/
test_input[7648:7655] = '{32'h41ac0cf8, 32'h41cf075b, 32'h42a67f33, 32'hc1214e10, 32'h416e9a87, 32'hc1c1ba37, 32'h41cb1d2d, 32'hc19fb58f};
test_label[956] = '{32'hc19fb58f};
test_output[956] = '{32'h42ce6c97};
/*############ DEBUG ############
test_input[7648:7655] = '{21.5063320814, 25.8785922349, 83.2484338921, -10.0815586601, 14.9127260466, -24.2159256791, 25.3892461884, -19.9636525358};
test_label[956] = '{-19.9636525358};
test_output[956] = '{103.212086428};
############ END DEBUG ############*/
test_input[7656:7663] = '{32'hc293f964, 32'h4279e72c, 32'hc282a43c, 32'hc23f1f29, 32'hc2c3080b, 32'h428dfdf0, 32'hc10ac869, 32'h41804ddc};
test_label[957] = '{32'hc293f964};
test_output[957] = '{32'h4310fbb7};
/*############ DEBUG ############
test_input[7656:7663] = '{-73.9870880465, 62.4757530846, -65.3207678569, -47.780430723, -97.5157122011, 70.99597157, -8.67392850021, 16.0380177246};
test_label[957] = '{-73.9870880465};
test_output[957] = '{144.983258992};
############ END DEBUG ############*/
test_input[7664:7671] = '{32'h426d4f8e, 32'hc24c807b, 32'hc2518736, 32'hc2368460, 32'hc26cf319, 32'hc265d226, 32'h412ca39f, 32'hc246e9ed};
test_label[958] = '{32'hc265d226};
test_output[958] = '{32'h42e990da};
/*############ DEBUG ############
test_input[7664:7671] = '{59.3276896783, -51.1254676166, -52.382041363, -45.6292713247, -59.2374011856, -57.4552231855, 10.7899464211, -49.7284439317};
test_label[958] = '{-57.4552231855};
test_output[958] = '{116.782912864};
############ END DEBUG ############*/
test_input[7672:7679] = '{32'hc2bb26c0, 32'hc1f4f45f, 32'h42b9d97a, 32'hc28a475e, 32'hc227925e, 32'hc1f50259, 32'hc28b6e42, 32'hc2c71d12};
test_label[959] = '{32'h42b9d97a};
test_output[959] = '{32'h80000000};
/*############ DEBUG ############
test_input[7672:7679] = '{-93.575684883, -30.6193209932, 92.9247557428, -69.1393905368, -41.8929381072, -30.6261457388, -69.7153445717, -99.5567817496};
test_label[959] = '{92.9247557428};
test_output[959] = '{-0.0};
############ END DEBUG ############*/
test_input[7680:7687] = '{32'hc17c7e61, 32'h414faf8e, 32'h41c52608, 32'h42460c94, 32'hc2042b4a, 32'hc1f27c6c, 32'hc0ec603a, 32'hc251aa48};
test_label[960] = '{32'h414faf8e};
test_output[960] = '{32'h421220b0};
/*############ DEBUG ############
test_input[7680:7687] = '{-15.7808544811, 12.9803604556, 24.6435696438, 49.5122822516, -33.0422732981, -30.3107524182, -7.38674633295, -52.4162898115};
test_label[960] = '{12.9803604556};
test_output[960] = '{36.531921796};
############ END DEBUG ############*/
test_input[7688:7695] = '{32'hc15d78e2, 32'h41819852, 32'h42054255, 32'h3fca979a, 32'h418a78e6, 32'hc12baffd, 32'hc2b80f11, 32'h42b66d80};
test_label[961] = '{32'hc15d78e2};
test_output[961] = '{32'h42d21c9c};
/*############ DEBUG ############
test_input[7688:7695] = '{-13.8420120618, 16.1993757228, 33.3147772717, 1.58275151292, 17.3090328847, -10.7304659673, -92.0294230002, 91.2138641206};
test_label[961] = '{-13.8420120618};
test_output[961] = '{105.055876182};
############ END DEBUG ############*/
test_input[7696:7703] = '{32'h42af74dc, 32'hc2bbba4c, 32'hc290764e, 32'h42a9ba12, 32'hc26e98c3, 32'hc1cac3d3, 32'h3f8d4a44, 32'hc2c793c2};
test_label[962] = '{32'hc2bbba4c};
test_output[962] = '{32'h4335a5c5};
/*############ DEBUG ############
test_input[7696:7703] = '{87.7282422189, -93.863864281, -72.2310646441, 84.86342091, -59.6491829735, -25.3456167082, 1.10382887453, -99.7885871598};
test_label[962] = '{-93.863864281};
test_output[962] = '{181.647534882};
############ END DEBUG ############*/
test_input[7704:7711] = '{32'h425a45ea, 32'hc26548aa, 32'hc20871b7, 32'hc24e49e5, 32'hc2ba5ba5, 32'hc291cbc7, 32'hc15f5c33, 32'hc292099c};
test_label[963] = '{32'h425a45ea};
test_output[963] = '{32'h80000000};
/*############ DEBUG ############
test_input[7704:7711] = '{54.5682743722, -57.3209604291, -34.1110494654, -51.5721621611, -93.1789928346, -72.8980024439, -13.9600092893, -73.0187712189};
test_label[963] = '{54.5682743722};
test_output[963] = '{-0.0};
############ END DEBUG ############*/
test_input[7712:7719] = '{32'hc28c4bb2, 32'hc1cc005a, 32'hc29cec99, 32'hc1ba93b2, 32'h4251bddf, 32'h428e2e8b, 32'hc2c21535, 32'hc283f753};
test_label[964] = '{32'h4251bddf};
test_output[964] = '{32'h41953e6e};
/*############ DEBUG ############
test_input[7712:7719] = '{-70.1478423096, -25.5001708915, -78.4621044347, -23.3221159157, 52.4354226767, 71.0909050662, -97.0414172972, -65.9830549048};
test_label[964] = '{52.4354226767};
test_output[964] = '{18.6554823974};
############ END DEBUG ############*/
test_input[7720:7727] = '{32'h42b53568, 32'h4221138f, 32'h41e22f9b, 32'hc2822d67, 32'hc1fc044f, 32'h42b8bd77, 32'h4210fc7e, 32'hc23cee5e};
test_label[965] = '{32'h42b8bd77};
test_output[965] = '{32'h3e21b30a};
/*############ DEBUG ############
test_input[7720:7727] = '{90.604305428, 40.2690990514, 28.2732442224, -65.0886727469, -31.5021042794, 92.3700448501, 36.2465762674, -47.2327811245};
test_label[965] = '{92.3700448501};
test_output[965] = '{0.157909538443};
############ END DEBUG ############*/
test_input[7728:7735] = '{32'h41e64eae, 32'h420de1b9, 32'h42c450dc, 32'h42bbbbc1, 32'hc2c16ba9, 32'h428ca9a6, 32'hc26c2563, 32'hc27b3b19};
test_label[966] = '{32'hc26c2563};
test_output[966] = '{32'h431d3542};
/*############ DEBUG ############
test_input[7728:7735] = '{28.788418436, 35.4704335754, 98.1579305675, 93.8667070065, -96.7102738658, 70.3313455137, -59.0365095633, -62.8077135818};
test_label[966] = '{-59.0365095633};
test_output[966] = '{157.208035461};
############ END DEBUG ############*/
test_input[7736:7743] = '{32'hc26cdc46, 32'hc1ed974c, 32'h428d3500, 32'hc28bfcd1, 32'hc2547068, 32'h40891db3, 32'h42437dca, 32'h41cb2480};
test_label[967] = '{32'h42437dca};
test_output[967] = '{32'h41add86e};
/*############ DEBUG ############
test_input[7736:7743] = '{-59.2151107958, -29.6988745736, 70.6035178028, -69.9937786381, -53.1097708601, 4.28487538888, 48.872839127, 25.3928224939};
test_label[967] = '{48.872839127};
test_output[967] = '{21.7306786762};
############ END DEBUG ############*/
test_input[7744:7751] = '{32'h42a934ee, 32'hc164b328, 32'h41f67f06, 32'hc2827bc5, 32'h428111ef, 32'h428caa0a, 32'h41d8a46e, 32'hc27c5fe3};
test_label[968] = '{32'h428111ef};
test_output[968] = '{32'h41a08bfb};
/*############ DEBUG ############
test_input[7744:7751] = '{84.6033780003, -14.2937396615, 30.812022238, -65.2417350175, 64.5350281631, 70.332104514, 27.0802878594, -63.0936396284};
test_label[968] = '{64.5350281631};
test_output[968] = '{20.0683504731};
############ END DEBUG ############*/
test_input[7752:7759] = '{32'hc0e33f51, 32'h4097b488, 32'hbfd6bb21, 32'h427bd331, 32'h417094f4, 32'h4232287f, 32'hc280d587, 32'hc1c779d6};
test_label[969] = '{32'hbfd6bb21};
test_output[969] = '{32'h42814485};
/*############ DEBUG ############
test_input[7752:7759] = '{-7.10147907207, 4.74078759941, -1.67758573528, 62.9562418321, 15.0363651533, 44.5395464913, -64.4170448866, -24.9344903991};
test_label[969] = '{-1.67758573528};
test_output[969] = '{64.6338275774};
############ END DEBUG ############*/
test_input[7760:7767] = '{32'h41bafa40, 32'h403990ca, 32'hc2ad8fd1, 32'hc29a2996, 32'h3f919600, 32'hc2b7d0f4, 32'h42ab3412, 32'h41952f7b};
test_label[970] = '{32'h41952f7b};
test_output[970] = '{32'h4285e833};
/*############ DEBUG ############
test_input[7760:7767] = '{23.3721916753, 2.89946211382, -86.7808900295, -77.0812234206, 1.1373901497, -91.9081097873, 85.6017003886, 18.6481844681};
test_label[970] = '{18.6481844681};
test_output[970] = '{66.9535159204};
############ END DEBUG ############*/
test_input[7768:7775] = '{32'hc276dbf1, 32'h42297c4a, 32'hc1c458df, 32'h41cb0037, 32'hc22ee9c8, 32'hc2a53e02, 32'hc275c37b, 32'hc1820bdc};
test_label[971] = '{32'hc275c37b};
test_output[971] = '{32'h42cf9fe3};
/*############ DEBUG ############
test_input[7768:7775] = '{-61.7147862174, 42.3713771351, -24.5433935671, 25.3751050135, -43.7283011833, -82.6211099959, -61.4408984771, -16.255790505};
test_label[971] = '{-61.4408984771};
test_output[971] = '{103.812275654};
############ END DEBUG ############*/
test_input[7776:7783] = '{32'h41e8840a, 32'h421a6865, 32'hc1e3b3c7, 32'hc1decd01, 32'h418867ff, 32'h42ab3703, 32'h427fe59b, 32'h41be84c7};
test_label[972] = '{32'hc1decd01};
test_output[972] = '{32'h42e2ea43};
/*############ DEBUG ############
test_input[7776:7783] = '{29.0644730421, 38.6019487073, -28.4627812692, -27.850100397, 17.0507798791, 85.6074444209, 63.9742251626, 23.8148327666};
test_label[972] = '{-27.850100397};
test_output[972] = '{113.457544818};
############ END DEBUG ############*/
test_input[7784:7791] = '{32'h41941389, 32'h42b0b7d9, 32'hc1e494eb, 32'hc178b657, 32'h41fda240, 32'hc296a5e3, 32'hc209a023, 32'h42bdcd45};
test_label[973] = '{32'hc296a5e3};
test_output[973] = '{32'h432a39f3};
/*############ DEBUG ############
test_input[7784:7791] = '{18.509538143, 88.3590763909, -28.5727146223, -15.5445164808, 31.7042240561, -75.3240008502, -34.406382853, 94.9009180028};
test_label[973] = '{-75.3240008502};
test_output[973] = '{170.226359645};
############ END DEBUG ############*/
test_input[7792:7799] = '{32'hc2a230cb, 32'h42ac09d5, 32'h3fab2480, 32'h41f09286, 32'h424e917f, 32'h4201b85a, 32'hc232ba77, 32'hc05c87f2};
test_label[974] = '{32'h3fab2480};
test_output[974] = '{32'h42a95d43};
/*############ DEBUG ############
test_input[7792:7799] = '{-81.0953024365, 86.0192040286, 1.33705140293, 30.0715442298, 51.642084362, 32.4300310248, -44.6820931014, -3.44579746846};
test_label[974] = '{1.33705140293};
test_output[974] = '{84.6821526257};
############ END DEBUG ############*/
test_input[7800:7807] = '{32'hc266f2c9, 32'h42c10778, 32'h4240e039, 32'h425512a6, 32'hc234a0a8, 32'h42c43216, 32'hc279e356, 32'h417a36be};
test_label[975] = '{32'h4240e039};
test_output[975] = '{32'h4248432c};
/*############ DEBUG ############
test_input[7800:7807] = '{-57.7370951253, 96.5145897972, 48.2189670084, 53.2682113158, -45.1568915386, 98.0978269356, -62.4720065566, 15.6383647768};
test_label[975] = '{48.2189670084};
test_output[975] = '{50.0655962299};
############ END DEBUG ############*/
test_input[7808:7815] = '{32'hc28c1749, 32'h4242027b, 32'h402394b9, 32'h41e669a4, 32'h4146d37b, 32'hc2a5d4ca, 32'hc25fa443, 32'h42018081};
test_label[976] = '{32'h4146d37b};
test_output[976] = '{32'h42104d9d};
/*############ DEBUG ############
test_input[7808:7815] = '{-70.0454756505, 48.5024231628, 2.55595231749, 28.8015825762, 12.4266305514, -82.9156049951, -55.9104134558, 32.3754903201};
test_label[976] = '{12.4266305514};
test_output[976] = '{36.0757927133};
############ END DEBUG ############*/
test_input[7816:7823] = '{32'h41802b2f, 32'hc2891703, 32'hc2a23d9b, 32'h42c7a9a5, 32'hc2afd7ac, 32'h41df3424, 32'h41e9d4ad, 32'hc2b5d61e};
test_label[977] = '{32'h41df3424};
test_output[977] = '{32'h428fdc9c};
/*############ DEBUG ############
test_input[7816:7823] = '{16.0210853142, -68.5449440276, -81.1203254305, 99.8313343473, -87.9212351129, 27.9004590251, 29.2288447255, -90.9182000029};
test_label[977] = '{27.9004590251};
test_output[977] = '{71.9308753223};
############ END DEBUG ############*/
test_input[7824:7831] = '{32'h41dd33d7, 32'h428f7bc1, 32'h42424cc6, 32'h42855743, 32'h420e0bfa, 32'h425724b2, 32'hc18cfabc, 32'hc136c825};
test_label[978] = '{32'h428f7bc1};
test_output[978] = '{32'h3bccf52d};
/*############ DEBUG ############
test_input[7824:7831] = '{27.6503129735, 71.7417099929, 48.5749755388, 66.6704324633, 35.5116943101, 53.7858341909, -17.6224294971, -11.423863156};
test_label[978] = '{71.7417099929};
test_output[978] = '{0.00625481310002};
############ END DEBUG ############*/
test_input[7832:7839] = '{32'h4212242b, 32'h42644f64, 32'h42614d9c, 32'h426f0aec, 32'h4212bf03, 32'h421e609f, 32'hc1ca8b3e, 32'h42293c02};
test_label[979] = '{32'h42614d9c};
test_output[979] = '{32'h4061f727};
/*############ DEBUG ############
test_input[7832:7839] = '{36.5353213108, 57.0775301445, 56.3257903147, 59.7606648166, 36.6865356979, 39.5943559922, -25.3179898686, 42.3086016841};
test_label[979] = '{56.3257903147};
test_output[979] = '{3.53071004426};
############ END DEBUG ############*/
test_input[7840:7847] = '{32'h427d455b, 32'h428338c1, 32'hc2bff1b3, 32'hc04528a3, 32'h42bccca3, 32'h41c54754, 32'h3ffafb4e, 32'hc0a50f68};
test_label[980] = '{32'h42bccca3};
test_output[980] = '{32'h2ac2c000};
/*############ DEBUG ############
test_input[7840:7847] = '{63.3177316267, 65.6108439914, -95.9720720002, -3.08060518906, 94.39967936, 24.6598290141, 1.96079425288, -5.15813065093};
test_label[980] = '{94.39967936};
test_output[980] = '{3.45945494473e-13};
############ END DEBUG ############*/
test_input[7848:7855] = '{32'h429e94a7, 32'hc1448200, 32'hc1834235, 32'h4069d92b, 32'h42097771, 32'h424ff579, 32'h42bbc4bb, 32'h42a78d6e};
test_label[981] = '{32'h429e94a7};
test_output[981] = '{32'h416980cc};
/*############ DEBUG ############
test_input[7848:7855] = '{79.2903369029, -12.2817379395, -16.4073269956, 3.65387988436, 34.3666429627, 51.9897185342, 93.8842399208, 83.7762317048};
test_label[981] = '{79.2903369029};
test_output[981] = '{14.5939442281};
############ END DEBUG ############*/
test_input[7856:7863] = '{32'hc233a0a6, 32'hc1088928, 32'h429565eb, 32'h42aa0b5c, 32'h40823efc, 32'h4209c44f, 32'hc2b63b6b, 32'hc24ad061};
test_label[982] = '{32'h429565eb};
test_output[982] = '{32'h41252baa};
/*############ DEBUG ############
test_input[7856:7863] = '{-44.9068839728, -8.53348509513, 74.6990590293, 85.0221867894, 4.07018842961, 34.4417073812, -91.1160510922, -50.7034958609};
test_label[982] = '{74.6990590293};
test_output[982] = '{10.3231606238};
############ END DEBUG ############*/
test_input[7864:7871] = '{32'h427ff711, 32'hc240ff42, 32'h41bce5eb, 32'h42180131, 32'h428c5e56, 32'h405fe02b, 32'hc13e3d03, 32'hc2172b7c};
test_label[983] = '{32'hc2172b7c};
test_output[983] = '{32'h42d7f51f};
/*############ DEBUG ############
test_input[7864:7871] = '{63.9912765981, -48.2492748573, 23.6122638924, 38.0011651887, 70.1842487021, 3.49805718655, -11.8898957943, -37.7924635634};
test_label[983] = '{-37.7924635634};
test_output[983] = '{107.978753923};
############ END DEBUG ############*/
test_input[7872:7879] = '{32'hc18386aa, 32'hc1bbc4f2, 32'h42b86770, 32'hc2a8098c, 32'hc1e82c2a, 32'hc2bf9d2a, 32'hc20a34c2, 32'hc2097bcb};
test_label[984] = '{32'hc18386aa};
test_output[984] = '{32'h42d9491a};
/*############ DEBUG ############
test_input[7872:7879] = '{-16.4407533229, -23.4711655307, 92.2020254907, -84.0186449032, -29.0215638277, -95.8069630951, -34.5515209303, -34.3708909077};
test_label[984] = '{-16.4407533229};
test_output[984] = '{108.642778814};
############ END DEBUG ############*/
test_input[7880:7887] = '{32'h429e910a, 32'hc27bc615, 32'h420af18d, 32'h4147bce1, 32'hc20ed387, 32'hc2bc662d, 32'hc0671a82, 32'hc2ab7517};
test_label[985] = '{32'h420af18d};
test_output[985] = '{32'h42323088};
/*############ DEBUG ############
test_input[7880:7887] = '{79.2832797008, -62.9434403414, 34.7358877194, 12.4836130274, -35.7065693187, -94.1995622303, -3.6109928753, -85.7286913539};
test_label[985] = '{34.7358877194};
test_output[985] = '{44.5473919814};
############ END DEBUG ############*/
test_input[7888:7895] = '{32'h42c583ab, 32'hc0ec7863, 32'hc29924a1, 32'h428a3f15, 32'hc1090b28, 32'h425a1ff9, 32'h42818b7f, 32'hc2bb9491};
test_label[986] = '{32'hc1090b28};
test_output[986] = '{32'h42d6a510};
/*############ DEBUG ############
test_input[7888:7895] = '{98.7571640355, -7.38969556351, -76.5715406949, 69.1232076808, -8.56522406201, 54.5312216969, 64.772452262, -93.7901655357};
test_label[986] = '{-8.56522406201};
test_output[986] = '{107.322388098};
############ END DEBUG ############*/
test_input[7896:7903] = '{32'h426884c8, 32'h41acdf81, 32'hc1a5aa88, 32'h40d9e703, 32'h41ac7d7e, 32'hc29d8163, 32'h42b6d232, 32'hc2a737b4};
test_label[987] = '{32'hc2a737b4};
test_output[987] = '{32'h432f04f3};
/*############ DEBUG ############
test_input[7896:7903] = '{58.1296706297, 21.6091336838, -20.7082672999, 6.80944975304, 21.5612762714, -78.7527105214, 91.4105365907, -83.6087947201};
test_label[987] = '{-83.6087947201};
test_output[987] = '{175.019331311};
############ END DEBUG ############*/
test_input[7904:7911] = '{32'h4168f866, 32'h42887fb0, 32'h421b61b8, 32'hc2ae01cf, 32'h423f5381, 32'h42671b73, 32'h4121c44d, 32'hc1ede793};
test_label[988] = '{32'h423f5381};
test_output[988] = '{32'h41a357cf};
/*############ DEBUG ############
test_input[7904:7911] = '{14.5606437504, 68.2493924789, 38.845428725, -87.0035311072, 47.8315458487, 57.7768071838, 10.1104250884, -29.7380732754};
test_label[988] = '{47.8315458487};
test_output[988] = '{20.4178749329};
############ END DEBUG ############*/
test_input[7912:7919] = '{32'h42735ebb, 32'h41b48e53, 32'h428d7c73, 32'hc28c5b50, 32'h3fdab147, 32'hc05dc043, 32'hc2c7e397, 32'hc1f3e047};
test_label[989] = '{32'hc05dc043};
test_output[989] = '{32'h42946a7c};
/*############ DEBUG ############
test_input[7912:7919] = '{60.8425084011, 22.5694938924, 70.7430647126, -70.1783439404, 1.70853506007, -3.46485963563, -99.9445134059, -30.4845097671};
test_label[989] = '{-3.46485963563};
test_output[989] = '{74.2079744938};
############ END DEBUG ############*/
test_input[7920:7927] = '{32'h4141c4c7, 32'hbe35ae16, 32'hc09f46f7, 32'h40df0dae, 32'h423105ad, 32'h41a0731b, 32'h427c5fa5, 32'hc297bd83};
test_label[990] = '{32'hc09f46f7};
test_output[990] = '{32'h42882442};
/*############ DEBUG ############
test_input[7920:7927] = '{12.110541495, -0.177421898565, -4.97741252487, 6.97041991019, 44.2555440579, 20.0562036884, 63.0934033621, -75.8701420644};
test_label[990] = '{-4.97741252487};
test_output[990] = '{68.0708158936};
############ END DEBUG ############*/
test_input[7928:7935] = '{32'hc27221a7, 32'hc269145a, 32'hc1f79dd1, 32'h42292838, 32'h42684d7f, 32'h4287a469, 32'h41bdacb2, 32'hc22cb7ff};
test_label[991] = '{32'hc269145a};
test_output[991] = '{32'h42fc2e9e};
/*############ DEBUG ############
test_input[7928:7935] = '{-60.5328636527, -58.269876347, -30.952058153, 42.2892754704, 58.0756787083, 67.8211164701, 23.7093230182, -43.179684888};
test_label[991] = '{-58.269876347};
test_output[991] = '{126.091051377};
############ END DEBUG ############*/
test_input[7936:7943] = '{32'h4255a2bc, 32'hc1a493db, 32'h41cbe0d4, 32'hc2619b80, 32'h42a9886a, 32'h4232fd50, 32'h4257bf6a, 32'hbfb1bb0c};
test_label[992] = '{32'hc1a493db};
test_output[992] = '{32'h42d2ad61};
/*############ DEBUG ############
test_input[7936:7943] = '{53.4089206104, -20.5721942871, 25.4847793212, -56.401855266, 84.7664331778, 44.7473773044, 53.9369270567, -1.3885207591};
test_label[992] = '{-20.5721942871};
test_output[992] = '{105.338627465};
############ END DEBUG ############*/
test_input[7944:7951] = '{32'hc2b7c036, 32'h42533c1e, 32'h42b6c182, 32'hc2ac35b8, 32'hbfb9027e, 32'hc2c2c6c0, 32'h40409f0a, 32'h42719a66};
test_label[993] = '{32'hc2b7c036};
test_output[993] = '{32'h433740dc};
/*############ DEBUG ############
test_input[7944:7951] = '{-91.8754158004, 52.8087074008, 91.3779424593, -86.1049231424, -1.44538857968, -97.3881852711, 3.00970689802, 60.4007814186};
test_label[993] = '{-91.8754158004};
test_output[993] = '{183.25335826};
############ END DEBUG ############*/
test_input[7952:7959] = '{32'hc2b0a979, 32'hc07000c9, 32'h41cd496a, 32'h429e82cc, 32'h4226c7de, 32'h4245cba0, 32'h423a3ab0, 32'h4151ca7f};
test_label[994] = '{32'hc2b0a979};
test_output[994] = '{32'h43279622};
/*############ DEBUG ############
test_input[7952:7959] = '{-88.3310038661, -3.7500479213, 25.66084639, 79.2554594649, 41.695180992, 49.4488536162, 46.5573114116, 13.1119372392};
test_label[994] = '{-88.3310038661};
test_output[994] = '{167.586463331};
############ END DEBUG ############*/
test_input[7960:7967] = '{32'h42a66ba4, 32'h421d70c3, 32'hc2775e9a, 32'hc21be328, 32'hc29f8c99, 32'h412d8b4b, 32'h421eccac, 32'h4127cc7e};
test_label[995] = '{32'hc21be328};
test_output[995] = '{32'h42f45d37};
/*############ DEBUG ############
test_input[7960:7967] = '{83.2102330887, 39.3601188515, -61.8423851226, -38.9718307915, -79.7746014531, 10.846507535, 39.699875351, 10.4874246507};
test_label[995] = '{-38.9718307915};
test_output[995] = '{122.18206388};
############ END DEBUG ############*/
test_input[7968:7975] = '{32'h42aeb632, 32'h428a327a, 32'hc1b85ecc, 32'hc101e7c2, 32'hc2baa8df, 32'hc24d72b0, 32'hc1cd7960, 32'h40a213c5};
test_label[996] = '{32'hc24d72b0};
test_output[996] = '{32'h430ab7c5};
/*############ DEBUG ############
test_input[7968:7975] = '{87.3558529854, 69.0985852992, -23.0462869758, -8.11908140015, -93.3298267593, -51.3619989953, -25.6842655383, 5.06491326481};
test_label[996] = '{-51.3619989953};
test_output[996] = '{138.717851992};
############ END DEBUG ############*/
test_input[7976:7983] = '{32'hc1fa8769, 32'hc2acefb4, 32'hc2b68ebb, 32'h42394afe, 32'h4299df19, 32'h429ad0ae, 32'h4193746f, 32'h41f5f54f};
test_label[997] = '{32'hc2acefb4};
test_output[997] = '{32'h43245c4d};
/*############ DEBUG ############
test_input[7976:7983] = '{-31.3161186642, -86.4681712322, -91.2787699271, 46.3232357495, 76.9357371683, 77.4075798326, 18.4318520689, 30.7447794607};
test_label[997] = '{-86.4681712322};
test_output[997] = '{164.36055196};
############ END DEBUG ############*/
test_input[7984:7991] = '{32'h429ef7aa, 32'hc2b34d14, 32'h420f5619, 32'h420f6c74, 32'h3da230c5, 32'hc2594f54, 32'h4215a773, 32'h42c58a34};
test_label[998] = '{32'hc2594f54};
test_output[998] = '{32'h431918ef};
/*############ DEBUG ############
test_input[7984:7991] = '{79.4837219103, -89.6505423361, 35.8340788426, 35.8559112973, 0.0791945795829, -54.3274695426, 37.413523295, 98.7699269731};
test_label[998] = '{-54.3274695426};
test_output[998] = '{153.09739652};
############ END DEBUG ############*/
test_input[7992:7999] = '{32'h41073c1f, 32'hc25db6c4, 32'h42b78cb3, 32'hc29149f8, 32'hc29a3fa7, 32'hc19ce17a, 32'h42bb9437, 32'hc29e8e56};
test_label[999] = '{32'h41073c1f};
test_output[999] = '{32'h42aaeccc};
/*############ DEBUG ############
test_input[7992:7999] = '{8.4521776839, -55.4284806292, 91.7748048065, -72.6444682472, -77.1243177142, -19.6100958049, 93.789478867, -79.27800109};
test_label[999] = '{8.4521776839};
test_output[999] = '{85.4624912652};
############ END DEBUG ############*/
test_input[8000:8007] = '{32'hc22fd178, 32'hc288a660, 32'h42c1d766, 32'hc260d9dc, 32'h419d8aa7, 32'hc21e754c, 32'h41413a9f, 32'hc1397588};
test_label[1000] = '{32'hc21e754c};
test_output[1000] = '{32'h43088906};
/*############ DEBUG ############
test_input[8000:8007] = '{-43.9545578825, -68.3249504975, 96.9207036945, -56.2127544105, 19.6927008598, -39.6145477641, 12.0768121479, -11.5911942827};
test_label[1000] = '{-39.6145477641};
test_output[1000] = '{136.535251459};
############ END DEBUG ############*/
test_input[8008:8015] = '{32'hc269530f, 32'hc28a8c78, 32'h429ddd8b, 32'h4062c56c, 32'hc202ecf6, 32'h40fee155, 32'hc2896aa2, 32'h42896664};
test_label[1001] = '{32'hc28a8c78};
test_output[1001] = '{32'h43143504};
/*############ DEBUG ############
test_input[8008:8015] = '{-58.3311119039, -69.2743520717, 78.9326973737, 3.54329963098, -32.7314078689, 7.96500647066, -68.708270543, 68.6999823473};
test_label[1001] = '{-69.2743520717};
test_output[1001] = '{148.207085419};
############ END DEBUG ############*/
test_input[8016:8023] = '{32'h42bc92d1, 32'hc1bf1c53, 32'hc203feca, 32'h425109c0, 32'h42877748, 32'h41e0d498, 32'h41a482ab, 32'hc239f3cb};
test_label[1002] = '{32'hc1bf1c53};
test_output[1002] = '{32'h42ec59e6};
/*############ DEBUG ############
test_input[8016:8023] = '{94.2867534963, -23.8888304698, -32.9988189273, 52.2595207196, 67.732970678, 28.1038050973, 20.5638019914, -46.4880801763};
test_label[1002] = '{-23.8888304698};
test_output[1002] = '{118.175583966};
############ END DEBUG ############*/
test_input[8024:8031] = '{32'hc2b9aa8c, 32'hc2ae3b9a, 32'hc288c212, 32'h42ae2451, 32'h42c1a300, 32'hc12d957b, 32'h41a96217, 32'h422785db};
test_label[1003] = '{32'hc2b9aa8c};
test_output[1003] = '{32'h433da6ca};
/*############ DEBUG ############
test_input[8024:8031] = '{-92.8330996762, -87.1164119925, -68.3790459166, 87.0709267715, 96.8183564274, -10.84899444, 21.1728960112, 41.8807176513};
test_label[1003] = '{-92.8330996762};
test_output[1003] = '{189.651514547};
############ END DEBUG ############*/
test_input[8032:8039] = '{32'h4284601e, 32'hc2a52d22, 32'h42033a21, 32'hbe56d6c5, 32'h42aa551f, 32'hc2c27c77, 32'h42be8b34, 32'hc1ed21f4};
test_label[1004] = '{32'hc2a52d22};
test_output[1004] = '{32'h4331dc2d};
/*############ DEBUG ############
test_input[8032:8039] = '{66.1877297552, -82.5881487964, 32.8067650394, -0.209803652405, 85.1662546656, -97.2430952665, 95.2718776213, -29.6415793552};
test_label[1004] = '{-82.5881487964};
test_output[1004] = '{177.860067266};
############ END DEBUG ############*/
test_input[8040:8047] = '{32'h41f7411a, 32'h41995574, 32'h4011a547, 32'hc296c2d4, 32'h4193b860, 32'hc2a321dd, 32'h4252b040, 32'h424bae98};
test_label[1005] = '{32'h4193b860};
test_output[1005] = '{32'h420977e3};
/*############ DEBUG ############
test_input[8040:8047] = '{30.9067869228, 19.1667248052, 2.27571279876, -75.3805210133, 18.4650273947, -81.5661377759, 52.6721186531, 50.920501658};
test_label[1005] = '{18.4650273947};
test_output[1005] = '{34.3670761824};
############ END DEBUG ############*/
test_input[8048:8055] = '{32'h42c4ea03, 32'h42ab16ce, 32'h41fb279a, 32'hc12a4631, 32'h423964c8, 32'hbf85dd70, 32'hc1236d11, 32'h425521bb};
test_label[1006] = '{32'h42c4ea03};
test_output[1006] = '{32'h36258e3f};
/*############ DEBUG ############
test_input[8048:8055] = '{98.457056965, 85.5445388874, 31.3943363884, -10.642136325, 46.3484186504, -1.04582025253, -10.214127256, 53.2829409367};
test_label[1006] = '{98.457056965};
test_output[1006] = '{2.46697140601e-06};
############ END DEBUG ############*/
test_input[8056:8063] = '{32'hc26d5c14, 32'hc2924272, 32'h41b104fd, 32'hc29b036a, 32'h42c23778, 32'h414f688a, 32'hc293e2ad, 32'hc2b8ddc0};
test_label[1007] = '{32'hc293e2ad};
test_output[1007] = '{32'h432b0d13};
/*############ DEBUG ############
test_input[8056:8063] = '{-59.3399182225, -73.1297733188, 22.1274364327, -77.5066704878, 97.1083352916, 12.9630224006, -73.9427285686, -92.4331029441};
test_label[1007] = '{-73.9427285686};
test_output[1007] = '{171.05106386};
############ END DEBUG ############*/
test_input[8064:8071] = '{32'h40b12d42, 32'h41837591, 32'h42b0b758, 32'h42006f3e, 32'hc1be52ed, 32'h41195f18, 32'hc273e51f, 32'hc1959fdb};
test_label[1008] = '{32'hc1959fdb};
test_output[1008] = '{32'h42d61f4f};
/*############ DEBUG ############
test_input[8064:8071] = '{5.53677443942, 16.4324058804, 88.3580968296, 32.1086338142, -23.7904916732, 9.58571667517, -60.9737524698, -18.7030539654};
test_label[1008] = '{-18.7030539654};
test_output[1008] = '{107.061150795};
############ END DEBUG ############*/
test_input[8072:8079] = '{32'hc27b9e0a, 32'h42b77fbf, 32'hc2a4538a, 32'h40d69768, 32'h42807383, 32'hc1b18a2d, 32'hc22a6bdb, 32'hc253a268};
test_label[1009] = '{32'hc253a268};
test_output[1009] = '{32'h4310a879};
/*############ DEBUG ############
test_input[8072:8079] = '{-62.904334437, 91.7495002884, -82.1631598046, 6.70598243172, 64.2256081756, -22.192468907, -42.6053283644, -52.908599863};
test_label[1009] = '{-52.908599863};
test_output[1009] = '{144.658100151};
############ END DEBUG ############*/
test_input[8080:8087] = '{32'hc29465d7, 32'h4253cf30, 32'hc2343346, 32'h42866db2, 32'hc219d5de, 32'h41748041, 32'hc29cf227, 32'hc28da7ee};
test_label[1010] = '{32'hc219d5de};
test_output[1010] = '{32'h42d358a1};
/*############ DEBUG ############
test_input[8080:8087] = '{-74.1989036548, 52.9523302435, -45.0500721306, 67.214252103, -38.4588542823, 15.28131226, -78.4729519877, -70.8279904597};
test_label[1010] = '{-38.4588542823};
test_output[1010] = '{105.673107025};
############ END DEBUG ############*/
test_input[8088:8095] = '{32'h4215f5ff, 32'hc2b41068, 32'hc29945ef, 32'h4288c60a, 32'h3fe8337a, 32'hc28dc188, 32'h3f8b132e, 32'hc11d014a};
test_label[1011] = '{32'h3fe8337a};
test_output[1011] = '{32'h4285253c};
/*############ DEBUG ############
test_input[8088:8095] = '{37.4902318446, -90.032042027, -76.6365895925, 68.38679563, 1.81407097209, -70.8779890955, 1.08652281042, -9.81281517472};
test_label[1011] = '{1.81407097209};
test_output[1011] = '{66.572724658};
############ END DEBUG ############*/
test_input[8096:8103] = '{32'h42982d61, 32'hc174f6a6, 32'hc1c41001, 32'h428742a8, 32'hc1f675d0, 32'h429afd15, 32'hc2024cdf, 32'h428d2123};
test_label[1012] = '{32'h428742a8};
test_output[1012] = '{32'h41215907};
/*############ DEBUG ############
test_input[8096:8103] = '{76.0886318216, -15.3102170671, -24.5078142451, 67.6301916425, -30.8075257673, 77.494300649, -32.5750698767, 70.5647168342};
test_label[1012] = '{67.6301916425};
test_output[1012] = '{10.0842347442};
############ END DEBUG ############*/
test_input[8104:8111] = '{32'h41aba5b3, 32'hc2c0e529, 32'h40d6a303, 32'hc2b03e4a, 32'h429b0c78, 32'h42c01349, 32'h42880518, 32'hc2975d13};
test_label[1013] = '{32'h429b0c78};
test_output[1013] = '{32'h41941b43};
/*############ DEBUG ############
test_input[8104:8111] = '{21.4559073292, -96.4475809387, 6.70739911572, -88.1216611923, 77.5243525729, 96.0376645455, 68.0099493847, -75.6817829259};
test_label[1013] = '{77.5243525729};
test_output[1013] = '{18.5133119817};
############ END DEBUG ############*/
test_input[8112:8119] = '{32'h42377969, 32'h424ef8cf, 32'hc284559f, 32'h424b3f7f, 32'hc1388631, 32'hc29cddbb, 32'h42c0bfb7, 32'hc083f2e8};
test_label[1014] = '{32'hc29cddbb};
test_output[1014] = '{32'h432eceb9};
/*############ DEBUG ############
test_input[8112:8119] = '{45.868564967, 51.7429760671, -66.1672318955, 50.8120073544, -11.532761248, -78.433070268, 96.3744442462, -4.12340187621};
test_label[1014] = '{-78.433070268};
test_output[1014] = '{174.807514514};
############ END DEBUG ############*/
test_input[8120:8127] = '{32'h4290e056, 32'h42b872e0, 32'hbf8ee9bd, 32'hc29e1343, 32'hc1891130, 32'h4147c187, 32'h42b32fcd, 32'hc192ae24};
test_label[1015] = '{32'hc192ae24};
test_output[1015] = '{32'h42dd4203};
/*############ DEBUG ############
test_input[8120:8127] = '{72.4381561984, 92.224365603, -1.11650809885, -79.0376199982, -17.1333920084, 12.4847482675, 89.5933627214, -18.3350299733};
test_label[1015] = '{-18.3350299733};
test_output[1015] = '{110.628927436};
############ END DEBUG ############*/
test_input[8128:8135] = '{32'h41a9fa01, 32'h42bb81b4, 32'h4230fc08, 32'hc1939d35, 32'h4288571b, 32'hc299de91, 32'hc2095528, 32'hc180f9e6};
test_label[1016] = '{32'hc1939d35};
test_output[1016] = '{32'h42e06901};
/*############ DEBUG ############
test_input[8128:8135] = '{21.2470722952, 93.753326962, 44.24612432, -18.4517617159, 68.1701291908, -76.9346988527, -34.3331605222, -16.1220207525};
test_label[1016] = '{-18.4517617159};
test_output[1016] = '{112.205088678};
############ END DEBUG ############*/
test_input[8136:8143] = '{32'hc1442315, 32'hc29e4d4c, 32'h4212e957, 32'hc28d6dba, 32'hc273de1f, 32'hc0fe49ff, 32'h41a7abbe, 32'hc2378a41};
test_label[1017] = '{32'hc29e4d4c};
test_output[1017] = '{32'h42e7c1f7};
/*############ DEBUG ############
test_input[8136:8143] = '{-12.2585651993, -79.1509696976, 36.7278705997, -70.7143072494, -60.9669151804, -7.94653264626, 20.9588588506, -45.8850146262};
test_label[1017] = '{-79.1509696976};
test_output[1017] = '{115.878840439};
############ END DEBUG ############*/
test_input[8144:8151] = '{32'h4248ef12, 32'h418d4004, 32'h42407a8c, 32'h42a53e81, 32'hc1c0e5de, 32'hc233342a, 32'h41e071bd, 32'h426f1e1c};
test_label[1018] = '{32'h41e071bd};
test_output[1018] = '{32'h425a4423};
/*############ DEBUG ############
test_input[8144:8151] = '{50.2334672089, 17.6562573543, 48.1196757377, 82.6220752866, -24.1122396568, -44.8009431103, 28.0555354859, 59.7794022209};
test_label[1018] = '{28.0555354859};
test_output[1018] = '{54.5665398008};
############ END DEBUG ############*/
test_input[8152:8159] = '{32'hc217c40f, 32'hc2a8df60, 32'h41c32656, 32'h423ab34a, 32'hc1d5cbf1, 32'h42a9ffcd, 32'h4281a901, 32'h422289e1};
test_label[1019] = '{32'hc2a8df60};
test_output[1019] = '{32'h43296f97};
/*############ DEBUG ############
test_input[8152:8159] = '{-37.9414623344, -84.4362770639, 24.3937196186, 46.6750862352, -26.7245810827, 84.9996132827, 64.8300884451, 40.6346483801};
test_label[1019] = '{-84.4362770639};
test_output[1019] = '{169.435890348};
############ END DEBUG ############*/
test_input[8160:8167] = '{32'hc2abda16, 32'h42a69656, 32'h41df5932, 32'hc166d07c, 32'h409caf01, 32'h423f3a18, 32'h427b9af3, 32'hc295f88d};
test_label[1020] = '{32'hc166d07c};
test_output[1020] = '{32'h42c37066};
/*############ DEBUG ############
test_input[8160:8167] = '{-85.9259514946, 83.2936257069, 27.9185531573, -14.4258994754, 4.89636279464, 47.8067339004, 62.9013190015, -74.9854505899};
test_label[1020] = '{-14.4258994754};
test_output[1020] = '{97.7195251837};
############ END DEBUG ############*/
test_input[8168:8175] = '{32'h42912a0b, 32'h428f3718, 32'h41724b5b, 32'h429438e5, 32'hc28cc4b7, 32'hc195ba58, 32'h42094123, 32'h41d71560};
test_label[1021] = '{32'h42912a0b};
test_output[1021] = '{32'h3fe5270c};
/*############ DEBUG ############
test_input[8168:8175] = '{72.5821114631, 71.6076076392, 15.1433973748, 74.1111188882, -70.3842107089, -18.7159885075, 34.3136088839, 26.8854373931};
test_label[1021] = '{72.5821114631};
test_output[1021] = '{1.79025413077};
############ END DEBUG ############*/
test_input[8176:8183] = '{32'hc20fa667, 32'hc2c00b20, 32'hc192dde1, 32'h418affb0, 32'hc28a794f, 32'h420a030a, 32'h42b70ccb, 32'h42156b72};
test_label[1022] = '{32'h420a030a};
test_output[1022] = '{32'h4264168d};
/*############ DEBUG ############
test_input[8176:8183] = '{-35.912501654, -96.0217320506, -18.3583395513, 17.3748479623, -69.2369286258, 34.5029661798, 91.5249891131, 37.3549255551};
test_label[1022] = '{34.5029661798};
test_output[1022] = '{57.0220229333};
############ END DEBUG ############*/
test_input[8184:8191] = '{32'hc235a7a4, 32'hc2326540, 32'hc1e037fc, 32'hc2ad9b31, 32'hc286fee6, 32'h40eff8a2, 32'h426ddd0c, 32'hc26adc86};
test_label[1023] = '{32'hc2326540};
test_output[1023] = '{32'h42d02126};
/*############ DEBUG ############
test_input[8184:8191] = '{-45.4137128387, -44.5988777526, -28.0273368041, -86.8031098652, -67.4978491239, 7.49910053584, 59.4658647048, -58.7153550404};
test_label[1023] = '{-44.5988777526};
test_output[1023] = '{104.064742457};
############ END DEBUG ############*/
test_input[8192:8199] = '{32'hc27a8aaa, 32'hc16245cd, 32'h41232096, 32'hc29185e2, 32'h42681d2d, 32'hc20c4995, 32'h4273d246, 32'h41f2da02};
test_label[1024] = '{32'h41232096};
test_output[1024] = '{32'h424b3f8f};
/*############ DEBUG ############
test_input[8192:8199] = '{-62.6354155176, -14.1420412559, 10.1954551743, -72.7614911225, 58.0284921012, -35.0718570945, 60.9553444946, 30.3564488083};
test_label[1024] = '{10.1954551743};
test_output[1024] = '{50.8120693284};
############ END DEBUG ############*/
test_input[8200:8207] = '{32'hc27a372c, 32'h42a08dc7, 32'hc2066a3a, 32'h42bea458, 32'hc2af942f, 32'h423d25fd, 32'hc290a024, 32'hc1f8f711};
test_label[1025] = '{32'hc2066a3a};
test_output[1025] = '{32'h4300ecbb};
/*############ DEBUG ############
test_input[8200:8207] = '{-62.5538791621, 80.2769070011, -33.6037363981, 95.3209862688, -87.789419853, 47.287096537, -72.3127775964, -31.1206383121};
test_label[1025] = '{-33.6037363981};
test_output[1025] = '{128.92472296};
############ END DEBUG ############*/
test_input[8208:8215] = '{32'h420bce9b, 32'hc16d738d, 32'hc29ed6ca, 32'hc2466ddb, 32'hc2117551, 32'hc1d63118, 32'hc2665a29, 32'h41cd1ae6};
test_label[1026] = '{32'hc2117551};
test_output[1026] = '{32'h428ea202};
/*############ DEBUG ############
test_input[8208:8215] = '{34.9517640551, -14.840710396, -79.4195088967, -49.6072798306, -36.3645659736, -26.7739720035, -57.5880480978, 25.638133893};
test_label[1026] = '{-36.3645659736};
test_output[1026] = '{71.3164202112};
############ END DEBUG ############*/
test_input[8216:8223] = '{32'h413db9e3, 32'hc20ab104, 32'hc0583610, 32'h429bf7d4, 32'h41b9113f, 32'h42b591d1, 32'hc23745f5, 32'hc2a1750b};
test_label[1027] = '{32'h42b591d1};
test_output[1027] = '{32'h3639219a};
/*############ DEBUG ############
test_input[8216:8223] = '{11.8578828799, -34.6728649951, -3.37829964893, 77.9840374596, 23.133421154, 90.7847977287, -45.8183183379, -80.7285959204};
test_label[1027] = '{90.7847977287};
test_output[1027] = '{2.75867063454e-06};
############ END DEBUG ############*/
test_input[8224:8231] = '{32'h42640b29, 32'hc2583a66, 32'hc28dd80c, 32'hbe876694, 32'h429ed09e, 32'h42c60c23, 32'h42526b17, 32'h4261a812};
test_label[1028] = '{32'hc28dd80c};
test_output[1028] = '{32'h4329f218};
/*############ DEBUG ############
test_input[8224:8231] = '{57.0108996925, -54.057029943, -70.9219683563, -0.264454493196, 79.4074577531, 99.0237043892, 52.604581016, 56.4141302491};
test_label[1028] = '{-70.9219683563};
test_output[1028] = '{169.945672749};
############ END DEBUG ############*/
test_input[8232:8239] = '{32'hc2138eb5, 32'h425905ef, 32'hc2b7c9e2, 32'h42b8a66a, 32'hc2597226, 32'hc2c6c66a, 32'hc2932949, 32'hc2b84a37};
test_label[1029] = '{32'hc2b7c9e2};
test_output[1029] = '{32'h43383826};
/*############ DEBUG ############
test_input[8232:8239] = '{-36.8893641566, 54.2557943029, -91.8943002765, 92.3250268966, -54.3614749179, -99.3875261565, -73.5806381566, -92.1449499974};
test_label[1029] = '{-91.8943002765};
test_output[1029] = '{184.219327173};
############ END DEBUG ############*/
test_input[8240:8247] = '{32'hc0650cab, 32'h427d099c, 32'h42c3e6ad, 32'hc27bf3a1, 32'h42a0ea63, 32'hc20fd01f, 32'hc1d48ec8, 32'h422de094};
test_label[1030] = '{32'hc0650cab};
test_output[1030] = '{32'h42cb0f12};
/*############ DEBUG ############
test_input[8240:8247] = '{-3.57889819587, 63.2593845484, 97.950534943, -62.9879177284, 80.4577842358, -35.9532418155, -26.5697172973, 43.4693153788};
test_label[1030] = '{-3.57889819587};
test_output[1030] = '{101.529433164};
############ END DEBUG ############*/
test_input[8248:8255] = '{32'hc1821e91, 32'h41a05a27, 32'hc292f62f, 32'hc2990c81, 32'hc298b1ee, 32'hc24f42bc, 32'hc2c6f6a5, 32'h42b81ddc};
test_label[1031] = '{32'h41a05a27};
test_output[1031] = '{32'h42900752};
/*############ DEBUG ############
test_input[8248:8255] = '{-16.264925114, 20.0440204956, -73.4808256146, -76.5244186656, -76.347519978, -51.8151701174, -99.4817293253, 92.0583186605};
test_label[1031] = '{20.0440204956};
test_output[1031] = '{72.014298165};
############ END DEBUG ############*/
test_input[8256:8263] = '{32'h42981ad6, 32'h424ebc9d, 32'h428a6417, 32'h42030417, 32'h42c09704, 32'hc16a15e5, 32'hc13ff61e, 32'hc224d017};
test_label[1032] = '{32'hc16a15e5};
test_output[1032] = '{32'h42ddd9c1};
/*############ DEBUG ############
test_input[8256:8263] = '{76.0524114733, 51.6841913682, 69.1954869481, 32.7539949321, 96.2949553808, -14.6303454317, -11.9975869237, -41.2032109091};
test_label[1032] = '{-14.6303454317};
test_output[1032] = '{110.925300814};
############ END DEBUG ############*/
test_input[8264:8271] = '{32'hc274764d, 32'hc254b6e6, 32'hc242aa4f, 32'h429149be, 32'h4256f2c7, 32'hc21a0a99, 32'hc047bebf, 32'hc29e2bdf};
test_label[1033] = '{32'hc21a0a99};
test_output[1033] = '{32'h42de4f0b};
/*############ DEBUG ############
test_input[8264:8271] = '{-61.1155277452, -53.1786126938, -48.6663187063, 72.6440292246, 53.7370885688, -38.5103486637, -3.12101718059, -79.0856863953};
test_label[1033] = '{-38.5103486637};
test_output[1033] = '{111.154377894};
############ END DEBUG ############*/
test_input[8272:8279] = '{32'hc2b6a3ab, 32'h428ae290, 32'hc2470f6e, 32'hc182b94c, 32'h41fb818e, 32'h42583b05, 32'h4279bdb5, 32'hc21c6930};
test_label[1034] = '{32'hc2470f6e};
test_output[1034] = '{32'h42ee6abe};
/*############ DEBUG ############
test_input[8272:8279] = '{-91.3196622151, 69.442508651, -49.7650695736, -16.3404775408, 31.4382594667, 54.0576373327, 62.4352602802, -39.1027239357};
test_label[1034] = '{-49.7650695736};
test_output[1034] = '{119.208483319};
############ END DEBUG ############*/
test_input[8280:8287] = '{32'hc2b55ed3, 32'hc29eb29d, 32'h4211f431, 32'hc211ecaf, 32'hc2707826, 32'h41051d49, 32'hc284675b, 32'hc1908a36};
test_label[1035] = '{32'hc2b55ed3};
test_output[1035] = '{32'h42fe58eb};
/*############ DEBUG ############
test_input[8280:8287] = '{-90.6852005909, -79.3488516965, 36.4884668454, -36.4811360482, -60.1173325815, 8.31964923483, -66.2018645074, -18.0674851466};
test_label[1035] = '{-90.6852005909};
test_output[1035] = '{127.173667436};
############ END DEBUG ############*/
test_input[8288:8295] = '{32'h4142e953, 32'h40634d33, 32'h415e55dd, 32'hc19aa32b, 32'h40be936e, 32'hc1e4d4cc, 32'h42c1bca1, 32'h42b9eb28};
test_label[1036] = '{32'h4142e953};
test_output[1036] = '{32'h42a969a2};
/*############ DEBUG ############
test_input[8288:8295] = '{12.1819635941, 3.55158686362, 13.8959624214, -19.3296727022, 5.95549655473, -28.6039055815, 96.868415546, 92.959289338};
test_label[1036] = '{12.1819635941};
test_output[1036] = '{84.7063114599};
############ END DEBUG ############*/
test_input[8296:8303] = '{32'hc2b254a4, 32'hc2c14e79, 32'h3fbba70c, 32'hc192c9af, 32'h42188676, 32'h42bae574, 32'h4282d39f, 32'h4176f6a0};
test_label[1037] = '{32'h4282d39f};
test_output[1037] = '{32'h41e04754};
/*############ DEBUG ############
test_input[8296:8303] = '{-89.165310887, -96.6532681681, 1.46603536663, -18.348479132, 38.1313079001, 93.4481491058, 65.4133205494, 15.4352111197};
test_label[1037] = '{65.4133205494};
test_output[1037] = '{28.0348285563};
############ END DEBUG ############*/
test_input[8304:8311] = '{32'h425fe8e0, 32'h422717c1, 32'h42a40567, 32'h42988b20, 32'hc20b119f, 32'h42a37eb5, 32'h4287734e, 32'hc28cedde};
test_label[1038] = '{32'h4287734e};
test_output[1038] = '{32'h416db7ec};
/*############ DEBUG ############
test_input[8304:8311] = '{55.9774170173, 41.7731957737, 82.0105501349, 76.2717289728, -34.7672072848, 81.747476248, 67.7252019563, -70.46458333};
test_label[1038] = '{67.7252019563};
test_output[1038] = '{14.857403014};
############ END DEBUG ############*/
test_input[8312:8319] = '{32'hc13cce67, 32'hc28ba63d, 32'h42401d77, 32'hc2a4d651, 32'hc0dffbb4, 32'h428dbaf2, 32'h4235632a, 32'hc09f9549};
test_label[1039] = '{32'hc28ba63d};
test_output[1039] = '{32'h430cb097};
/*############ DEBUG ############
test_input[8312:8319] = '{-11.8003913973, -69.824683262, 48.0287756984, -82.4185851167, -6.99947566255, 70.8651281571, 45.3468383753, -4.98697332221};
test_label[1039] = '{-69.824683262};
test_output[1039] = '{140.689811419};
############ END DEBUG ############*/
test_input[8320:8327] = '{32'hc14af205, 32'h42b96610, 32'hc12fa87b, 32'h418a802c, 32'hc2833e25, 32'hc1f4308e, 32'h42a00064, 32'hc29347e1};
test_label[1040] = '{32'hc29347e1};
test_output[1040] = '{32'h432656f9};
/*############ DEBUG ############
test_input[8320:8327] = '{-12.684086504, 92.699340483, -10.9786329703, 17.3125848635, -65.621375191, -30.5237091732, 80.0007649547, -73.6403886561};
test_label[1040] = '{-73.6403886561};
test_output[1040] = '{166.339732195};
############ END DEBUG ############*/
test_input[8328:8335] = '{32'hc1579310, 32'hc29ca878, 32'h41c231a8, 32'h42937775, 32'h424708dc, 32'hc2957501, 32'hc26460ce, 32'hc22177de};
test_label[1041] = '{32'h424708dc};
test_output[1041] = '{32'h41bfcc1d};
/*############ DEBUG ############
test_input[8328:8335] = '{-13.473404349, -78.3290422352, 24.2742455884, 73.7333152667, 49.7586503993, -74.7285225259, -57.0945375178, -40.3670567954};
test_label[1041] = '{49.7586503993};
test_output[1041] = '{23.9746648675};
############ END DEBUG ############*/
test_input[8336:8343] = '{32'h42bb10d1, 32'h41ce39be, 32'h42a3461e, 32'h42301420, 32'hc23cf36b, 32'h4291691a, 32'h4145478a, 32'hc24e270c};
test_label[1042] = '{32'h42301420};
test_output[1042] = '{32'h42460d84};
/*############ DEBUG ############
test_input[8336:8343] = '{93.5328465007, 25.7781944791, 81.6369439509, 44.0196551869, -47.2377145595, 72.7052745316, 12.3299655216, -51.5381307126};
test_label[1042] = '{44.0196551869};
test_output[1042] = '{49.513198133};
############ END DEBUG ############*/
test_input[8344:8351] = '{32'hc2bb0a98, 32'h40b96b67, 32'h42693f47, 32'h41a2cfde, 32'hc2ac24dd, 32'hc2ab0cbf, 32'h4227499a, 32'hc27bc29b};
test_label[1043] = '{32'h41a2cfde};
test_output[1043] = '{32'h4217d758};
/*############ DEBUG ############
test_input[8344:8351] = '{-93.5206930229, 5.79436074267, 58.3117950645, 20.3514982374, -86.0719975891, -85.5248979684, 41.821877973, -62.9400461505};
test_label[1043] = '{20.3514982374};
test_output[1043] = '{37.960296896};
############ END DEBUG ############*/
test_input[8352:8359] = '{32'h40b45cc8, 32'hc29daa0a, 32'hc2ac5349, 32'hc12dce43, 32'hc246f897, 32'h429d3066, 32'hc1d14543, 32'hc196392f};
test_label[1044] = '{32'hc29daa0a};
test_output[1044] = '{32'h431d6d38};
/*############ DEBUG ############
test_input[8352:8359] = '{5.63632561109, -78.8321108019, -86.1626678208, -10.8628572995, -49.7427618867, 78.5945247567, -26.1588198694, -18.7779223586};
test_label[1044] = '{-78.8321108019};
test_output[1044] = '{157.426635559};
############ END DEBUG ############*/
test_input[8360:8367] = '{32'hc1e8b8f1, 32'hc2bd6b4c, 32'hc197c335, 32'hc2550a39, 32'h42ad4fea, 32'hc255922b, 32'h420ac0f6, 32'hc277047f};
test_label[1045] = '{32'hc255922b};
test_output[1045] = '{32'h430c0c80};
/*############ DEBUG ############
test_input[8360:8367] = '{-29.0903034015, -94.7095672787, -18.9703166174, -53.259983451, 86.6560800739, -53.3927418031, 34.6884395665, -61.7543917924};
test_label[1045] = '{-53.3927418031};
test_output[1045] = '{140.048821877};
############ END DEBUG ############*/
test_input[8368:8375] = '{32'hc1ab934f, 32'h412644ce, 32'hc2a59900, 32'h422c49a9, 32'hc2057a60, 32'hc2a2a50c, 32'hc14e8cbc, 32'h429b477e};
test_label[1046] = '{32'h412644ce};
test_output[1046] = '{32'h42867ee5};
/*############ DEBUG ############
test_input[8368:8375] = '{-21.4469288453, 10.3917978794, -82.7988312891, 43.0719335573, -33.3695066215, -81.322357252, -12.9093592166, 77.639635212};
test_label[1046] = '{10.3917978794};
test_output[1046] = '{67.2478373326};
############ END DEBUG ############*/
test_input[8376:8383] = '{32'h42c1deed, 32'h42133357, 32'h4150a83d, 32'h41029d82, 32'hc08c2b90, 32'hc27057e7, 32'h4086e312, 32'hc2a13608};
test_label[1047] = '{32'hc27057e7};
test_output[1047] = '{32'h431d0570};
/*############ DEBUG ############
test_input[8376:8383] = '{96.9354015448, 36.8001363758, 13.0410739824, 8.16345452717, -4.38031788519, -60.0858407782, 4.2152187041, -80.6055283952};
test_label[1047] = '{-60.0858407782};
test_output[1047] = '{157.021242323};
############ END DEBUG ############*/
test_input[8384:8391] = '{32'h42aa3c47, 32'hc2026dee, 32'hc1ce8b9a, 32'hc1a4e090, 32'hc2c20cd6, 32'hc0179577, 32'h417c7041, 32'hc282360c};
test_label[1048] = '{32'hc2026dee};
test_output[1048] = '{32'h42eb733e};
/*############ DEBUG ############
test_input[8384:8391] = '{85.1177263918, -32.6073537218, -25.8181646144, -20.6096503201, -97.0250685995, -2.36849770429, 15.7774054387, -65.105556914};
test_label[1048] = '{-32.6073537218};
test_output[1048] = '{117.725080114};
############ END DEBUG ############*/
test_input[8392:8399] = '{32'h42b3b96b, 32'hc1920e77, 32'hc1ddc3e6, 32'h421813c9, 32'hc25ed665, 32'h42b1c6be, 32'h422e40f2, 32'hc27f9c19};
test_label[1049] = '{32'h42b3b96b};
test_output[1049] = '{32'h3ea401fe};
/*############ DEBUG ############
test_input[8392:8399] = '{89.8621438287, -18.2570634034, -27.7206539168, 38.0193222371, -55.7093706481, 88.888168709, 43.5634224952, -63.9024379393};
test_label[1049] = '{89.8621438287};
test_output[1049] = '{0.320327704131};
############ END DEBUG ############*/
test_input[8400:8407] = '{32'h4299c33a, 32'h42aeca6c, 32'h428c4d9a, 32'h4283c651, 32'h42af6115, 32'hc2a4919c, 32'h4270a36d, 32'hc1ffefa3};
test_label[1050] = '{32'h42aeca6c};
test_output[1050] = '{32'h3f59dfd9};
/*############ DEBUG ############
test_input[8400:8407] = '{76.8813015207, 87.3953532443, 70.1515674767, 65.8873357147, 87.6896103158, -82.2843959888, 60.1595970856, -31.9920100754};
test_label[1050] = '{87.3953532443};
test_output[1050] = '{0.85107190157};
############ END DEBUG ############*/
test_input[8408:8415] = '{32'hc2a7448d, 32'h3f9ff550, 32'h41bc2887, 32'hc212da9b, 32'h42b09510, 32'hc22995f8, 32'h4210963a, 32'hc21c9534};
test_label[1051] = '{32'hc212da9b};
test_output[1051] = '{32'h42fa025d};
/*############ DEBUG ############
test_input[8408:8415] = '{-83.6338893481, 1.24967387285, 23.5197884689, -36.7134814641, 88.2911360905, -42.3964547735, 36.1467037929, -39.1457050363};
test_label[1051] = '{-36.7134814641};
test_output[1051] = '{125.004617555};
############ END DEBUG ############*/
test_input[8416:8423] = '{32'hc2500867, 32'h429670d5, 32'h427b6c3e, 32'h41330604, 32'h42b6a28d, 32'h410f01ce, 32'hc282e4ad, 32'hc24ea31d};
test_label[1052] = '{32'h42b6a28d};
test_output[1052] = '{32'h33db4dd2};
/*############ DEBUG ############
test_input[8416:8423] = '{-52.0082065406, 75.220373414, 62.8557046194, 11.1889683301, 91.3174813881, 8.93794053794, -65.4466295849, -51.659290444};
test_label[1052] = '{91.3174813881};
test_output[1052] = '{1.02121377129e-07};
############ END DEBUG ############*/
test_input[8424:8431] = '{32'hc27d4021, 32'hc1f151d3, 32'h4134ac27, 32'hc1a85ef1, 32'hc29c3b2c, 32'hc1f2fbb0, 32'hc088a298, 32'hc23f368a};
test_label[1053] = '{32'hc1f2fbb0};
test_output[1053] = '{32'h4226a8e2};
/*############ DEBUG ############
test_input[8424:8431] = '{-63.3126276599, -30.1649533197, 11.2920290218, -21.046357929, -78.115571166, -30.3728944521, -4.26984783276, -47.8032608127};
test_label[1053] = '{-30.3728944521};
test_output[1053] = '{41.6649236483};
############ END DEBUG ############*/
test_input[8432:8439] = '{32'hc028b402, 32'hc16f274b, 32'h418524bd, 32'hc2aa9490, 32'hc1b88479, 32'hc299c3da, 32'hc284e24f, 32'hc216f90c};
test_label[1054] = '{32'h418524bd};
test_output[1054] = '{32'h3191a752};
/*############ DEBUG ############
test_input[8432:8439] = '{-2.63598689048, -14.94709322, 16.6429378371, -85.2901645882, -23.0646839802, -76.8825242191, -66.4420063764, -37.7432110979};
test_label[1054] = '{16.6429378371};
test_output[1054] = '{4.23907732038e-09};
############ END DEBUG ############*/
test_input[8440:8447] = '{32'h42884e62, 32'h424c5eae, 32'hc2b74db3, 32'hc2174625, 32'h41ad423c, 32'h419f5e40, 32'hc285fb3a, 32'h42ae666b};
test_label[1055] = '{32'h42884e62};
test_output[1055] = '{32'h41986022};
/*############ DEBUG ############
test_input[8440:8447] = '{68.1530939439, 51.092461488, -91.6517575266, -37.8185021327, 21.6573415074, 19.9210203837, -66.9906740989, 87.2000336946};
test_label[1055] = '{68.1530939439};
test_output[1055] = '{19.0469397561};
############ END DEBUG ############*/
test_input[8448:8455] = '{32'hc1da89b3, 32'h42ba8bac, 32'h404ecd1a, 32'hc2adbd42, 32'h427bfe07, 32'hc299fa0e, 32'hc0cf3a94, 32'hc27f5eec};
test_label[1056] = '{32'h404ecd1a};
test_output[1056] = '{32'h42b41543};
/*############ DEBUG ############
test_input[8448:8455] = '{-27.3172364691, 93.2727964947, 3.23126832029, -86.8696455173, 62.9980730398, -76.9883853423, -6.47590072855, -63.8426984158};
test_label[1056] = '{3.23126832029};
test_output[1056] = '{90.0415281744};
############ END DEBUG ############*/
test_input[8456:8463] = '{32'hc0e4cc41, 32'h4185ba17, 32'h429f2941, 32'hc24235c8, 32'hc184d018, 32'hc29ac5f5, 32'hc24c40fe, 32'hc2b61821};
test_label[1057] = '{32'h429f2941};
test_output[1057] = '{32'h80000000};
/*############ DEBUG ############
test_input[8456:8463] = '{-7.14993349878, 16.7158635322, 79.580575106, -48.5525198841, -16.6016084632, -77.3866356809, -51.0634691148, -91.0471296572};
test_label[1057] = '{79.580575106};
test_output[1057] = '{-0.0};
############ END DEBUG ############*/
test_input[8464:8471] = '{32'h420a9736, 32'h42c55000, 32'hc23ff988, 32'hc2894398, 32'h42b03d3d, 32'hc2a9beb2, 32'hc2a3fca5, 32'hc1ca31d1};
test_label[1058] = '{32'h42c55000};
test_output[1058] = '{32'h37deadb9};
/*############ DEBUG ############
test_input[8464:8471] = '{34.647665619, 98.6562515955, -47.9936842948, -68.6320199508, 88.1196091885, -84.8724501833, -81.9934440499, -25.2743249276};
test_label[1058] = '{98.6562515955};
test_output[1058] = '{2.65453576239e-05};
############ END DEBUG ############*/
test_input[8472:8479] = '{32'hc286d2be, 32'h422cd481, 32'h42434efb, 32'hc21c3b4c, 32'hc2837488, 32'h42b883b4, 32'h42c73d06, 32'h4299848f};
test_label[1059] = '{32'hc286d2be};
test_output[1059] = '{32'h4327080c};
/*############ DEBUG ############
test_input[8472:8479] = '{-67.4116076601, 43.2075245051, 48.8271297514, -39.0579087372, -65.7275972979, 92.2572335884, 99.6191875746, 76.7589070481};
test_label[1059] = '{-67.4116076601};
test_output[1059] = '{167.03142999};
############ END DEBUG ############*/
test_input[8480:8487] = '{32'h424eb4f3, 32'h41ef2e59, 32'hc1da1bf8, 32'hc285c1ab, 32'hc2a5a0eb, 32'h41031bcb, 32'h424f2ae3, 32'hc1afcd0c};
test_label[1060] = '{32'hc1da1bf8};
test_output[1060] = '{32'h429f62b1};
/*############ DEBUG ############
test_input[8480:8487] = '{51.6767067347, 29.897629826, -27.263657297, -66.8782542404, -82.8142929221, 8.19428529858, 51.7918810211, -21.9751201295};
test_label[1060] = '{-27.263657297};
test_output[1060] = '{79.6927555794};
############ END DEBUG ############*/
test_input[8488:8495] = '{32'h421db2e0, 32'hc2b56aa4, 32'h424561e0, 32'h425bc6b9, 32'hc22a4185, 32'h4230a9dc, 32'hc27ad472, 32'hc24e31b7};
test_label[1061] = '{32'hc27ad472};
test_output[1061] = '{32'h42eb4f7d};
/*############ DEBUG ############
test_input[8488:8495] = '{39.424683066, -90.7082854749, 49.3455803497, 54.944064289, -42.563984105, 44.1658781628, -62.7074677498, -51.5485509461};
test_label[1061] = '{-62.7074677498};
test_output[1061] = '{117.655249625};
############ END DEBUG ############*/
test_input[8496:8503] = '{32'h428253b2, 32'h4269c950, 32'hc2b0501d, 32'h424e4e2b, 32'h428933b2, 32'hc2035402, 32'hc0fc142a, 32'h421e9752};
test_label[1062] = '{32'h424e4e2b};
test_output[1062] = '{32'h41887351};
/*############ DEBUG ############
test_input[8496:8503] = '{65.1634707874, 58.4465953163, -88.156471814, 51.5763376587, 68.6009684733, -32.8320387589, -7.87746140451, 39.6477729382};
test_label[1062] = '{51.5763376587};
test_output[1062] = '{17.0563077291};
############ END DEBUG ############*/
test_input[8504:8511] = '{32'hc2ae8288, 32'hc2a0236c, 32'hc27ff8d1, 32'hc2a9d17d, 32'hc26ee9e1, 32'hc214a3c9, 32'h422e3b57, 32'hc2c02943};
test_label[1063] = '{32'hc2a9d17d};
test_output[1063] = '{32'h43007794};
/*############ DEBUG ############
test_input[8504:8511] = '{-87.2549413709, -80.0691814987, -63.9929830239, -84.9091567484, -59.7283985094, -37.1599452754, 43.5579474807, -96.0805887599};
test_label[1063] = '{-84.9091567484};
test_output[1063] = '{128.467104229};
############ END DEBUG ############*/
test_input[8512:8519] = '{32'h428c78bb, 32'hc2b05819, 32'hc2aedb75, 32'h42bdc752, 32'hc21f5672, 32'hc29b2f42, 32'h42b09dfc, 32'hc0cd1883};
test_label[1064] = '{32'h428c78bb};
test_output[1064] = '{32'h41c53d33};
/*############ DEBUG ############
test_input[8512:8519] = '{70.2358028695, -88.1720622363, -87.4286251267, 94.889300275, -39.8344182615, -77.5923023727, 88.3085641534, -6.4092421648};
test_label[1064] = '{70.2358028695};
test_output[1064] = '{24.6548832729};
############ END DEBUG ############*/
test_input[8520:8527] = '{32'hc2c7e347, 32'hc29ba5ae, 32'h42848779, 32'h42c6ccfd, 32'h41cde894, 32'h423f8229, 32'hc261e35c, 32'h42b460ec};
test_label[1065] = '{32'h42c6ccfd};
test_output[1065] = '{32'h38d18d56};
/*############ DEBUG ############
test_input[8520:8527] = '{-99.9438993975, -77.8235964244, 66.2645944406, 99.4003686431, 25.7385634789, 47.8771087851, -56.4720293821, 90.1893001783};
test_label[1065] = '{99.4003686431};
test_output[1065] = '{9.99222248294e-05};
############ END DEBUG ############*/
test_input[8528:8535] = '{32'h422ad361, 32'h42720e69, 32'hc2807a08, 32'hc2af8fd3, 32'h423c3ef8, 32'h429a2f85, 32'h40e9b302, 32'h42b2ae34};
test_label[1066] = '{32'hc2807a08};
test_output[1066] = '{32'h4319941e};
/*############ DEBUG ############
test_input[8528:8535] = '{42.7064251259, 60.5140734406, -64.2383413104, -87.7809056906, 47.0614937019, 77.0928113993, 7.30310176421, 89.3402400742};
test_label[1066] = '{-64.2383413104};
test_output[1066] = '{153.578586182};
############ END DEBUG ############*/
test_input[8536:8543] = '{32'hc2966d68, 32'h42a00310, 32'hc2405299, 32'hc2272b9c, 32'h4134c86d, 32'h4160bad6, 32'hc245b534, 32'hc1b2d7d2};
test_label[1067] = '{32'h42a00310};
test_output[1067] = '{32'h80000000};
/*############ DEBUG ############
test_input[8536:8543] = '{-75.2136825841, 80.0059826727, -48.0806606817, -41.7925881641, 11.2989317524, 14.0456145376, -49.4269549163, -22.3553817253};
test_label[1067] = '{80.0059826727};
test_output[1067] = '{-0.0};
############ END DEBUG ############*/
test_input[8544:8551] = '{32'h42260c75, 32'h42c6a2c9, 32'hc2c415f1, 32'hc2725bdf, 32'hc1648da9, 32'hc18615e9, 32'hc28e77d1, 32'hc20ed53d};
test_label[1068] = '{32'hc2725bdf};
test_output[1068] = '{32'h431fe85c};
/*############ DEBUG ############
test_input[8544:8551] = '{41.5121664985, 99.3179406145, -98.0428565132, -60.5897170231, -14.2845853675, -16.7606980818, -71.2340188109, -35.7082417143};
test_label[1068] = '{-60.5897170231};
test_output[1068] = '{159.907657638};
############ END DEBUG ############*/
test_input[8552:8559] = '{32'hc2a52503, 32'hc22676ee, 32'h41ec5106, 32'h42bf9d90, 32'h41d18605, 32'hc241ee57, 32'h428fbe5b, 32'hc2c3f114};
test_label[1069] = '{32'h428fbe5b};
test_output[1069] = '{32'h41bf7cd4};
/*############ DEBUG ############
test_input[8552:8559] = '{-82.5722878067, -41.6161410664, 29.539562136, 95.8077381856, 26.190440053, -48.4827548114, 71.8717874913, -97.9708590867};
test_label[1069] = '{71.8717874913};
test_output[1069] = '{23.9359506943};
############ END DEBUG ############*/
test_input[8560:8567] = '{32'hbf876caa, 32'h40c65a45, 32'h42a81375, 32'h42c60d51, 32'hc285deb9, 32'h42c4a99b, 32'hc2b66b0b, 32'hc1f68a9a};
test_label[1070] = '{32'h42a81375};
test_output[1070] = '{32'h41764976};
/*############ DEBUG ############
test_input[8560:8567] = '{-1.05800361999, 6.19851918759, 84.0380043133, 99.0260068094, -66.9350038738, 98.3312586983, -91.2090716711, -30.8176765128};
test_label[1070] = '{84.0380043133};
test_output[1070] = '{15.3929344519};
############ END DEBUG ############*/
test_input[8568:8575] = '{32'h420e8bbb, 32'hc2101af2, 32'hc049d940, 32'h42907ee7, 32'hc22e6139, 32'h41aea81f, 32'hc123902a, 32'h4255b134};
test_label[1071] = '{32'hc22e6139};
test_output[1071] = '{32'h42e7af84};
/*############ DEBUG ############
test_input[8568:8575] = '{35.6364563186, -36.0263122111, -3.15388479733, 72.2478559341, -43.5949456139, 21.8320894463, -10.2226965551, 53.4230484443};
test_label[1071] = '{-43.5949456139};
test_output[1071] = '{115.842801555};
############ END DEBUG ############*/
test_input[8576:8583] = '{32'hc2902018, 32'h429e7870, 32'h41a41176, 32'hc21cb203, 32'h413bf43b, 32'hc27f1414, 32'hc1c8e1c3, 32'h41944127};
test_label[1072] = '{32'h429e7870};
test_output[1072] = '{32'h80000000};
/*############ DEBUG ############
test_input[8576:8583] = '{-72.0626838764, 79.2352288222, 20.5085257117, -39.1738400236, 11.7471269568, -63.7696063459, -25.110236122, 18.5318125455};
test_label[1072] = '{79.2352288222};
test_output[1072] = '{-0.0};
############ END DEBUG ############*/
test_input[8584:8591] = '{32'h42c2da0c, 32'h41c24dd7, 32'hc1e4bad5, 32'h428c7bc4, 32'hc1ca3166, 32'h4201e54c, 32'h408431f4, 32'hc185024a};
test_label[1073] = '{32'hc1ca3166};
test_output[1073] = '{32'h42f56665};
/*############ DEBUG ############
test_input[8584:8591] = '{97.4258724906, 24.2880082345, -28.5912270078, 70.241726059, -25.2741198886, 32.4739223885, 4.13109784246, -16.6261170364};
test_label[1073] = '{-25.2741198886};
test_output[1073] = '{122.699992379};
############ END DEBUG ############*/
test_input[8592:8599] = '{32'hc269cb2f, 32'h42070b18, 32'h4280bb82, 32'h42a138f0, 32'hc2535712, 32'h4231aec1, 32'hc2a20ca9, 32'hc02b08d4};
test_label[1074] = '{32'hc02b08d4};
test_output[1074] = '{32'h42a69136};
/*############ DEBUG ############
test_input[8592:8599] = '{-58.4484223961, 33.7608347669, 64.3662241839, 80.6112048872, -52.8350303462, 44.4206584996, -81.0247276447, -2.67241391222};
test_label[1074] = '{-2.67241391222};
test_output[1074] = '{83.2836188875};
############ END DEBUG ############*/
test_input[8600:8607] = '{32'hc16524c1, 32'h4212d41e, 32'hc29e47a0, 32'h42c732fb, 32'h428b6027, 32'h42aa6cdb, 32'h42bedbac, 32'hc29f4145};
test_label[1075] = '{32'hc16524c1};
test_output[1075] = '{32'h42e3df6c};
/*############ DEBUG ############
test_input[8600:8607] = '{-14.3214730852, 36.7071460117, -79.1398894257, 99.5995713207, 69.6877956312, 85.2126066503, 95.4290429535, -79.6274822382};
test_label[1075] = '{-14.3214730852};
test_output[1075] = '{113.936371014};
############ END DEBUG ############*/
test_input[8608:8615] = '{32'hc2bbe390, 32'h41823d17, 32'h4141771b, 32'hc2a7ce04, 32'h4219df2e, 32'h42a7b066, 32'hc2a18ba0, 32'h402daa55};
test_label[1076] = '{32'h4141771b};
test_output[1076] = '{32'h428f8183};
/*############ DEBUG ############
test_input[8608:8615] = '{-93.9444616813, 16.2798287816, 12.0915785082, -83.9023715779, 38.4679501724, 83.8445299485, -80.7727076362, 2.71352133315};
test_label[1076] = '{12.0915785082};
test_output[1076] = '{71.7529514404};
############ END DEBUG ############*/
test_input[8616:8623] = '{32'h4156580d, 32'hc248f3f8, 32'hc228e695, 32'hc28b2747, 32'hc1a7120e, 32'hc132b612, 32'hc12e7f23, 32'hc2086319};
test_label[1077] = '{32'hc1a7120e};
test_output[1077] = '{32'h42091f0a};
/*############ DEBUG ############
test_input[8616:8623] = '{13.3964969497, -50.2382526319, -42.2251778552, -69.5767112975, -20.8838162075, -11.1694509751, -10.9060396469, -34.0967747452};
test_label[1077] = '{-20.8838162075};
test_output[1077] = '{34.2803131573};
############ END DEBUG ############*/
test_input[8624:8631] = '{32'hc1819d20, 32'hc231d90f, 32'h41d90b66, 32'h412cbff3, 32'hc2b25957, 32'h427c1166, 32'hc2aa0aa3, 32'h41d64b4c};
test_label[1078] = '{32'hc231d90f};
test_output[1078] = '{32'h42d6f53a};
/*############ DEBUG ############
test_input[8624:8631] = '{-16.2017211085, -44.461972386, 27.130566092, 10.7968622969, -89.1744907627, 63.0169887678, -85.020772234, 26.7867660899};
test_label[1078] = '{-44.461972386};
test_output[1078] = '{107.478961154};
############ END DEBUG ############*/
test_input[8632:8639] = '{32'hc2b354bb, 32'hc2bfe2aa, 32'hc2b18e7c, 32'h42747fce, 32'hc2c62f99, 32'hc13fe6f9, 32'h42a8cc8e, 32'hc1b5f2f4};
test_label[1079] = '{32'hc2b18e7c};
test_output[1079] = '{32'h432d2d85};
/*############ DEBUG ############
test_input[8632:8639] = '{-89.6654898062, -95.9427042163, -88.7782931235, 61.1248099366, -99.0929668166, -11.9938895863, 84.3995220228, -22.7436303588};
test_label[1079] = '{-88.7782931235};
test_output[1079] = '{173.177815146};
############ END DEBUG ############*/
test_input[8640:8647] = '{32'hc19f8a2f, 32'hc29534ad, 32'h420d052f, 32'h40a08b25, 32'h4258a2d4, 32'hc174ede6, 32'hc282ea38, 32'hc21bd35a};
test_label[1080] = '{32'h40a08b25};
test_output[1080] = '{32'h42449170};
/*############ DEBUG ############
test_input[8640:8647] = '{-19.9424727793, -74.6028856532, 35.2550603998, 5.01698553195, 54.159012887, -15.3080810935, -65.4574569406, -38.9563977471};
test_label[1080] = '{5.01698553195};
test_output[1080] = '{49.1420273612};
############ END DEBUG ############*/
test_input[8648:8655] = '{32'hc045963c, 32'hc2414c51, 32'h42ad3cc7, 32'h41cbcb4a, 32'h4244be45, 32'hc2590889, 32'hc294f582, 32'h40aa4f16};
test_label[1081] = '{32'hc294f582};
test_output[1081] = '{32'h43211924};
/*############ DEBUG ############
test_input[8648:8655] = '{-3.0872944836, -48.3245291629, 86.6187030249, 25.4742627274, 49.1858088339, -54.2583351243, -74.4795070982, 5.32215384029};
test_label[1081] = '{-74.4795070982};
test_output[1081] = '{161.098210123};
############ END DEBUG ############*/
test_input[8656:8663] = '{32'h42b58064, 32'hc28294f3, 32'h42b895a0, 32'hc2046c61, 32'hc2a4a919, 32'h421e42ab, 32'h42181a7c, 32'hc2a36d54};
test_label[1082] = '{32'hc2a36d54};
test_output[1082] = '{32'h432e3322};
/*############ DEBUG ############
test_input[8656:8663] = '{90.7507612782, -65.2909168207, 92.2922350941, -33.1058382377, -82.3302672494, 39.5651041892, 38.0258654899, -81.7135341052};
test_label[1082] = '{-81.7135341052};
test_output[1082] = '{174.199743742};
############ END DEBUG ############*/
test_input[8664:8671] = '{32'h42778188, 32'h42b129dc, 32'hc299988f, 32'hc25ce067, 32'h422f8d9b, 32'h4053f03a, 32'h41c46c8e, 32'hc2714805};
test_label[1083] = '{32'h42778188};
test_output[1083] = '{32'h41d5a45e};
/*############ DEBUG ############
test_input[8664:8671] = '{61.8764972234, 88.5817538065, -76.7979637343, -55.2191430573, 43.8882850525, 3.31153735872, 24.5530060709, -60.3203330664};
test_label[1083] = '{61.8764972234};
test_output[1083] = '{26.7052565831};
############ END DEBUG ############*/
test_input[8672:8679] = '{32'h419cab2b, 32'hc2a193f8, 32'h41927c1e, 32'hc2836680, 32'h425251a0, 32'h42b70101, 32'hc271273a, 32'hc29d6f18};
test_label[1084] = '{32'h425251a0};
test_output[1084] = '{32'h421bb062};
/*############ DEBUG ############
test_input[8672:8679] = '{19.5835785659, -80.7890051341, 18.3106036362, -65.7001964584, 52.5797112053, 91.5019584469, -60.2883055465, -78.7169776798};
test_label[1084] = '{52.5797112053};
test_output[1084] = '{38.9222472416};
############ END DEBUG ############*/
test_input[8680:8687] = '{32'h423b53f7, 32'h422a13ca, 32'hc2457328, 32'hc279e363, 32'hc28d81ce, 32'h428a2605, 32'hc1820b3f, 32'h42ac8173};
test_label[1085] = '{32'h42ac8173};
test_output[1085] = '{32'h3314bb1a};
/*############ DEBUG ############
test_input[8680:8687] = '{46.8319952492, 42.5193239812, -49.3624562806, -62.472056297, -70.7535273148, 69.0742606881, -16.2554917866, 86.2528320521};
test_label[1085] = '{86.2528320521};
test_output[1085] = '{3.4629102963e-08};
############ END DEBUG ############*/
test_input[8688:8695] = '{32'h425da34a, 32'hc2789738, 32'hc2ad993f, 32'hc250b654, 32'h4253bb69, 32'h41bbdc0a, 32'hc29a05ff, 32'hc238fa0f};
test_label[1086] = '{32'h41bbdc0a};
test_output[1086] = '{32'h420007e7};
/*############ DEBUG ############
test_input[8688:8695] = '{55.4094602038, -62.1476751327, -86.7993088113, -52.1780542468, 52.9330196331, 23.482441301, -77.0117126113, -46.2441976001};
test_label[1086] = '{23.482441301};
test_output[1086] = '{32.0077153981};
############ END DEBUG ############*/
test_input[8696:8703] = '{32'h427ec09b, 32'h429f8ebf, 32'h4210b7fa, 32'hc27b340a, 32'hc28f3477, 32'hc2bb3e6b, 32'hc1ea67ae, 32'hc2b8db85};
test_label[1087] = '{32'hc28f3477};
test_output[1087] = '{32'h4317619b};
/*############ DEBUG ############
test_input[8696:8703] = '{63.6880904867, 79.7788035186, 36.1796637918, -62.8008177026, -71.6024740153, -93.6219093762, -29.3006244899, -92.4287462764};
test_label[1087] = '{-71.6024740153};
test_output[1087] = '{151.381277637};
############ END DEBUG ############*/
test_input[8704:8711] = '{32'hc1ebf721, 32'h420c7e89, 32'hc2384661, 32'h424927af, 32'hc1398a7e, 32'h424e4c1d, 32'hc08fd523, 32'hc2ad115c};
test_label[1088] = '{32'hc1ebf721};
test_output[1088] = '{32'h42a2a0d3};
/*############ DEBUG ############
test_input[8704:8711] = '{-29.4956678297, 35.1235684406, -46.0687308289, 50.2887529789, -11.596311609, 51.5743276601, -4.49476757574, -86.5339068996};
test_label[1088] = '{-29.4956678297};
test_output[1088] = '{81.3141109572};
############ END DEBUG ############*/
test_input[8712:8719] = '{32'hc203848b, 32'h4224d8de, 32'h4115cb99, 32'hc2b0a775, 32'h4272fb8e, 32'hc2062d86, 32'h42a5b479, 32'hc26daa08};
test_label[1089] = '{32'h4115cb99};
test_output[1089] = '{32'h4292fb06};
/*############ DEBUG ############
test_input[8712:8719] = '{-32.8794371596, 41.2117846007, 9.36220658289, -88.3270626994, 60.7456589086, -33.5444577161, 82.8524829324, -59.4160474488};
test_label[1089] = '{9.36220658289};
test_output[1089] = '{73.4902763497};
############ END DEBUG ############*/
test_input[8720:8727] = '{32'h4241c50b, 32'h40e3a79b, 32'hc268f185, 32'hc26a6580, 32'h4276bfe3, 32'h4265d7bb, 32'hc2275a96, 32'h4195a2d5};
test_label[1090] = '{32'h40e3a79b};
test_output[1090] = '{32'h425a59c8};
/*############ DEBUG ############
test_input[8720:8727] = '{48.4424257606, 7.11420952151, -58.235859399, -58.5991206793, 61.6873892835, 57.4606756496, -41.8384643337, 18.7045075815};
test_label[1090] = '{7.11420952151};
test_output[1090] = '{54.5876762414};
############ END DEBUG ############*/
test_input[8728:8735] = '{32'h41812a5a, 32'h428098a4, 32'h428801be, 32'h40792ce1, 32'hc13e3320, 32'hc286eb23, 32'hc29d1a11, 32'h41dbab8b};
test_label[1091] = '{32'hc286eb23};
test_output[1091] = '{32'h43077ca9};
/*############ DEBUG ############
test_input[8728:8735] = '{16.1456794185, 64.2981295928, 68.0033991292, 3.8933641308, -11.8874812143, -67.4592540237, -78.5509120362, 27.4587612348};
test_label[1091] = '{-67.4592540237};
test_output[1091] = '{135.486949187};
############ END DEBUG ############*/
test_input[8736:8743] = '{32'h4296d4eb, 32'h42ae2859, 32'hc2b97d61, 32'h419e7ab0, 32'h4214fb96, 32'h41a6e716, 32'hc18b0060, 32'h429717ee};
test_label[1092] = '{32'h429717ee};
test_output[1092] = '{32'h41388365};
/*############ DEBUG ############
test_input[8736:8743] = '{75.4158578286, 87.0788005291, -92.7448823449, 19.8099066554, 37.2456894489, 20.8628355816, -17.3751829895, 75.5467405424};
test_label[1092] = '{75.5467405424};
test_output[1092] = '{11.5320784039};
############ END DEBUG ############*/
test_input[8744:8751] = '{32'hc185e250, 32'h42b31a31, 32'h419ff4a3, 32'hc0960241, 32'h429b19c9, 32'h425bfe62, 32'hc21af3e1, 32'hc184b690};
test_label[1093] = '{32'h425bfe62};
test_output[1093] = '{32'h420a3600};
/*############ DEBUG ############
test_input[8744:8751] = '{-16.7355046892, 89.5511522848, 19.9944516094, -4.68777495172, 77.55035794, 54.9984225216, -38.738161566, -16.5891418173};
test_label[1093] = '{54.9984225216};
test_output[1093] = '{34.5527359025};
############ END DEBUG ############*/
test_input[8752:8759] = '{32'h4184a35d, 32'h425994df, 32'h420769b5, 32'h429f3215, 32'hc2a1eae6, 32'h42777a8c, 32'h42ad195e, 32'hc145008d};
test_label[1094] = '{32'h425994df};
test_output[1094] = '{32'h42009ed7};
/*############ DEBUG ############
test_input[8752:8759] = '{16.5797680121, 54.3953811953, 33.8532314259, 79.5978165628, -80.9587832964, 61.869675703, 86.5495433032, -12.3126340722};
test_label[1094] = '{54.3953811953};
test_output[1094] = '{32.1551186315};
############ END DEBUG ############*/
test_input[8760:8767] = '{32'h41ffcace, 32'hc15b51a6, 32'h40abddd8, 32'h4274048e, 32'h4244a971, 32'h42b80788, 32'h423da691, 32'hc11c6058};
test_label[1095] = '{32'h4244a971};
test_output[1095] = '{32'h422b659e};
/*############ DEBUG ############
test_input[8760:8767] = '{31.9740255821, -13.7074332587, 5.37083060458, 61.0044484157, 49.1654696613, 92.0147070621, 47.4126633173, -9.77352112264};
test_label[1095] = '{49.1654696613};
test_output[1095] = '{42.8492374008};
############ END DEBUG ############*/
test_input[8768:8775] = '{32'h42c02ce8, 32'h42146557, 32'hc2916f68, 32'hc2a96f5a, 32'hc28dc8cc, 32'h4283f5ca, 32'h42b57192, 32'hc2bdef1c};
test_label[1096] = '{32'hc2a96f5a};
test_output[1096] = '{32'h4334cf53};
/*############ DEBUG ############
test_input[8768:8775] = '{96.0877097622, 37.0989659738, -72.7175869851, -84.7174870591, -70.8921795011, 65.9800538839, 90.7218136955, -94.9670123028};
test_label[1096] = '{-84.7174870591};
test_output[1096] = '{180.809859206};
############ END DEBUG ############*/
test_input[8776:8783] = '{32'hc2b6d168, 32'hc2a540af, 32'h422b2b6b, 32'hc2bf0433, 32'h425c9aa1, 32'h41b2feaf, 32'hc29ac9ec, 32'h414d22df};
test_label[1097] = '{32'h422b2b6b};
test_output[1097] = '{32'h4145bcdd};
/*############ DEBUG ############
test_input[8776:8783] = '{-91.4089932762, -82.6263386945, 42.7923985892, -95.5082030104, 55.1510036727, 22.3743576054, -77.3943775254, 12.8210132563};
test_label[1097] = '{42.7923985892};
test_output[1097] = '{12.3586093761};
############ END DEBUG ############*/
test_input[8784:8791] = '{32'h4188f5e3, 32'hc1ce929f, 32'h426e6d27, 32'hc29775f4, 32'h429eed1e, 32'h427ca736, 32'h418067da, 32'hc238422f};
test_label[1098] = '{32'h426e6d27};
test_output[1098] = '{32'h419eda2c};
/*############ DEBUG ############
test_input[8784:8791] = '{17.1200619887, -25.8215931606, 59.6065931884, -75.7303783395, 79.4631226882, 63.1632903898, 16.0507082188, -46.0646321471};
test_label[1098] = '{59.6065931884};
test_output[1098] = '{19.8565295856};
############ END DEBUG ############*/
test_input[8792:8799] = '{32'h40ce1e28, 32'h420cf456, 32'hc1420e1d, 32'h41a645ab, 32'h420ed4d3, 32'hc2c16594, 32'h41500684, 32'hc26f3448};
test_label[1099] = '{32'h41500684};
test_output[1099] = '{32'h41b98953};
/*############ DEBUG ############
test_input[8792:8799] = '{6.44118096475, 35.2386100894, -12.1284453696, 20.7840175008, 35.707837056, -96.6983976897, 13.0015903197, -59.8010570818};
test_label[1099] = '{13.0015903197};
test_output[1099] = '{23.1920535431};
############ END DEBUG ############*/
test_input[8800:8807] = '{32'h421aafe9, 32'h42a49395, 32'hc1086958, 32'h4084046e, 32'hc28dcb78, 32'hc2523381, 32'h40c813fe, 32'hc2b12472};
test_label[1100] = '{32'hc28dcb78};
test_output[1100] = '{32'h43192f87};
/*############ DEBUG ############
test_input[8800:8807] = '{38.6717864607, 82.2882466267, -8.52571845377, 4.12554089514, -70.89740112, -52.5502954557, 6.25244053633, -88.5711843617};
test_label[1100] = '{-70.89740112};
test_output[1100] = '{153.185647747};
############ END DEBUG ############*/
test_input[8808:8815] = '{32'h42c5965f, 32'h41540026, 32'h42ba6833, 32'h421405f9, 32'h4203c129, 32'h42904003, 32'hc16be52e, 32'hc2b3b901};
test_label[1101] = '{32'h41540026};
test_output[1101] = '{32'h42ab1843};
/*############ DEBUG ############
test_input[8808:8815] = '{98.7936957535, 13.2500358147, 93.2035157308, 37.0058311787, 32.9386327873, 72.1250244361, -14.7434521251, -89.8613336557};
test_label[1101] = '{13.2500358147};
test_output[1101] = '{85.5473873389};
############ END DEBUG ############*/
test_input[8816:8823] = '{32'h426c0442, 32'hc28b99f2, 32'h3f9e1c45, 32'h429aa4f3, 32'h41e684e6, 32'hc2b70504, 32'h41e0b874, 32'hc236cb8e};
test_label[1102] = '{32'h41e0b874};
test_output[1102] = '{32'h4244edab};
/*############ DEBUG ############
test_input[8816:8823] = '{59.0041593256, -69.8006743296, 1.23523769646, 77.3221640314, 28.8148916714, -91.5097977198, 28.0900648741, -45.6987820824};
test_label[1102] = '{28.0900648741};
test_output[1102] = '{49.2320991684};
############ END DEBUG ############*/
test_input[8824:8831] = '{32'h41af4c69, 32'hc28f8018, 32'hc115950a, 32'hc2c2ba23, 32'hc28095d1, 32'h418b98c4, 32'hc24610a8, 32'hc22c44ba};
test_label[1103] = '{32'hc2c2ba23};
test_output[1103] = '{32'h42ee931c};
/*############ DEBUG ############
test_input[8824:8831] = '{21.9123101015, -71.7501830906, -9.34888652937, -97.363548901, -64.2926083535, 17.4495933928, -49.516267613, -43.0671175439};
test_label[1103] = '{-97.363548901};
test_output[1103] = '{119.287324022};
############ END DEBUG ############*/
test_input[8832:8839] = '{32'hc2746e83, 32'hc2b0008d, 32'h4241fcbd, 32'h42166ec9, 32'h42c3810b, 32'h40c4e400, 32'hc28c33cf, 32'hc20b46eb};
test_label[1104] = '{32'h42c3810b};
test_output[1104] = '{32'h80000000};
/*############ DEBUG ############
test_input[8832:8839] = '{-61.1079223917, -88.0010778859, 48.4968149309, 37.6081880172, 97.7520397839, 6.15283205736, -70.1011868839, -34.8192546755};
test_label[1104] = '{97.7520397839};
test_output[1104] = '{-0.0};
############ END DEBUG ############*/
test_input[8840:8847] = '{32'h42b0bf9b, 32'h4184faca, 32'hc1ebb490, 32'hc28738c8, 32'hc2b649b5, 32'hc2a04dc2, 32'h41f067a2, 32'h42b68339};
test_label[1105] = '{32'hc1ebb490};
test_output[1105] = '{32'h42f18c45};
/*############ DEBUG ############
test_input[8840:8847] = '{88.3742265075, 16.6224552351, -29.4631661858, -67.6108999523, -91.1439579707, -80.1518691983, 30.0506026395, 91.2562926095};
test_label[1105] = '{-29.4631661858};
test_output[1105] = '{120.77396488};
############ END DEBUG ############*/
test_input[8848:8855] = '{32'h421fdf2f, 32'hc2a6d28d, 32'hc28557d7, 32'h4106efad, 32'hc2a9dead, 32'hc2b10fed, 32'h42029396, 32'h42ab4d59};
test_label[1106] = '{32'hc2a9dead};
test_output[1106] = '{32'h432a9603};
/*############ DEBUG ############
test_input[8848:8855] = '{39.9679537256, -83.4112325582, -66.6715645461, 8.43351468102, -84.934912335, -88.5311030755, 32.6441257952, 85.6510713503};
test_label[1106] = '{-84.934912335};
test_output[1106] = '{170.585983685};
############ END DEBUG ############*/
test_input[8856:8863] = '{32'h429fa350, 32'hc27e036c, 32'h41999dde, 32'hc10681e9, 32'hc2a0f4e2, 32'h42912c97, 32'h42a8113d, 32'hc23db8fa};
test_label[1107] = '{32'hc2a0f4e2};
test_output[1107] = '{32'h432486d2};
/*############ DEBUG ############
test_input[8856:8863] = '{79.8189696325, -63.50334254, 19.2020827478, -8.40671628008, -80.4782873538, 72.5870903811, 84.0336678938, -47.4306420702};
test_label[1107] = '{-80.4782873538};
test_output[1107] = '{164.526634445};
############ END DEBUG ############*/
test_input[8864:8871] = '{32'h42249af6, 32'hc28fb162, 32'h42c34d48, 32'h4297641a, 32'hbeef5975, 32'h426ad2e8, 32'hc23ce409, 32'h4232ae07};
test_label[1108] = '{32'hc23ce409};
test_output[1108] = '{32'h4310dfa6};
/*############ DEBUG ############
test_input[8864:8871] = '{41.1513283364, -71.8464511032, 97.6509365702, 75.6955073119, -0.467479367614, 58.7059634117, -47.2226890443, 44.669949075};
test_label[1108] = '{-47.2226890443};
test_output[1108] = '{144.873625615};
############ END DEBUG ############*/
test_input[8872:8879] = '{32'hc25c0cce, 32'hc28559bf, 32'h41b3919c, 32'h4268c4f4, 32'h41314098, 32'h4103aa8c, 32'hc1681251, 32'hc2c1e8fe};
test_label[1109] = '{32'h41b3919c};
test_output[1109] = '{32'h420efc26};
/*############ DEBUG ############
test_input[8872:8879] = '{-55.0125051917, -66.6752888145, 22.4460988973, 58.1923376, 11.0782703869, 8.22913728593, -14.5044716358, -96.9550594551};
test_label[1109] = '{22.4460988973};
test_output[1109] = '{35.7462387027};
############ END DEBUG ############*/
test_input[8880:8887] = '{32'h428162c1, 32'h42a8dc81, 32'hc2b7633a, 32'hbf8bca2f, 32'hc2aa12d2, 32'hc0c59dab, 32'h42395e48, 32'hc2828fa4};
test_label[1110] = '{32'hc2b7633a};
test_output[1110] = '{32'h43301fdd};
/*############ DEBUG ############
test_input[8880:8887] = '{64.6928772679, 84.4306706865, -91.6937982072, -1.09210766543, -85.0367567961, -6.1754967987, 46.3420730492, -65.2805461504};
test_label[1110] = '{-91.6937982072};
test_output[1110] = '{176.124468896};
############ END DEBUG ############*/
test_input[8888:8895] = '{32'h42310885, 32'h42819727, 32'h4280ea4f, 32'hbf8446b5, 32'hc1991a84, 32'hc2037c95, 32'h42ac3e3d, 32'hc2b3fbc3};
test_label[1111] = '{32'hc1991a84};
test_output[1111] = '{32'h42d284de};
/*############ DEBUG ############
test_input[8888:8895] = '{44.2583208399, 64.7952224486, 64.4576326213, -1.03340778579, -19.1379476765, -32.8716615308, 86.1215557511, -89.9917233251};
test_label[1111] = '{-19.1379476765};
test_output[1111] = '{105.259503429};
############ END DEBUG ############*/
test_input[8896:8903] = '{32'hc1cf3af7, 32'hc265e852, 32'h4172b4f7, 32'h42a4fb3a, 32'hc2124aaa, 32'hc2b86f2e, 32'h413ddd85, 32'hc115b6b9};
test_label[1112] = '{32'hc265e852};
test_output[1112] = '{32'h430bf7b2};
/*############ DEBUG ############
test_input[8896:8903] = '{-25.9037907605, -57.4768771419, 15.1691812521, 82.4906765048, -36.572914034, -92.2171466389, 11.8665823748, -9.35711005297};
test_label[1112] = '{-57.4768771419};
test_output[1112] = '{139.967553647};
############ END DEBUG ############*/
test_input[8904:8911] = '{32'h42843dd1, 32'hc216d250, 32'h41297391, 32'hc297bec3, 32'hc261fe64, 32'hc2b95a97, 32'h41bbfdcb, 32'h41df687e};
test_label[1113] = '{32'h41df687e};
test_output[1113] = '{32'h4218c763};
/*############ DEBUG ############
test_input[8904:8911] = '{66.1207342513, -37.7053846055, 10.5907140809, -75.8725777077, -56.4984264777, -92.6769359435, 23.4989220132, 27.9260219872};
test_label[1113] = '{27.9260219872};
test_output[1113] = '{38.1947122641};
############ END DEBUG ############*/
test_input[8912:8919] = '{32'h42afa848, 32'hc28bb3ba, 32'hc1fee28a, 32'hc2a08283, 32'h42923e95, 32'h42b42cc8, 32'h42ab6855, 32'h425cc899};
test_label[1114] = '{32'h42923e95};
test_output[1114] = '{32'h41889b52};
/*############ DEBUG ############
test_input[8912:8919] = '{87.828676206, -69.8510281719, -31.8606142239, -80.2549054821, 73.1222310939, 90.087464082, 85.7037768917, 55.1958957592};
test_label[1114] = '{73.1222310939};
test_output[1114] = '{17.0758404298};
############ END DEBUG ############*/
test_input[8920:8927] = '{32'hc2824a1d, 32'h4292b78b, 32'h4267b7b9, 32'hc283936e, 32'h42bcc211, 32'hc23351fb, 32'h42aba816, 32'hc1d10f6a};
test_label[1115] = '{32'h42aba816};
test_output[1115] = '{32'h4108d0a0};
/*############ DEBUG ############
test_input[8920:8927] = '{-65.1447523035, 73.3584823927, 57.9294157756, -65.7879458671, 94.3790362883, -44.8300577808, 85.8282960815, -26.1325262241};
test_label[1115] = '{85.8282960815};
test_output[1115] = '{8.55093359073};
############ END DEBUG ############*/
test_input[8928:8935] = '{32'h429a41c0, 32'h40a2b078, 32'h428d2ba4, 32'hc1ddaea3, 32'h42427aa9, 32'hc28c3498, 32'h42654eb7, 32'hc1fa0508};
test_label[1116] = '{32'h428d2ba4};
test_output[1116] = '{32'h40d16d86};
/*############ DEBUG ############
test_input[8928:8935] = '{77.1284196803, 5.08404176767, 70.5852390974, -27.7102711696, 48.6197852457, -70.1027195327, 57.3268693682, -31.2524573202};
test_label[1116] = '{70.5852390974};
test_output[1116] = '{6.54461945125};
############ END DEBUG ############*/
test_input[8936:8943] = '{32'h427203b7, 32'hc2a1a746, 32'hc292ee13, 32'hc2bb5ed3, 32'h41f51f8d, 32'hc1fdaace, 32'hc2c2e0d2, 32'hc0d101b5};
test_label[1117] = '{32'hc2a1a746};
test_output[1117] = '{32'h430d5491};
/*############ DEBUG ############
test_input[8936:8943] = '{60.5036271208, -80.8267092625, -73.4649918439, -93.6852003226, 30.6404064898, -31.7084014372, -97.4391022333, -6.53145860373};
test_label[1117] = '{-80.8267092625};
test_output[1117] = '{141.330336383};
############ END DEBUG ############*/
test_input[8944:8951] = '{32'hc2201c66, 32'hc2c4b36e, 32'hc1b7d1b7, 32'hc1d20978, 32'hc21e8cb3, 32'h42c4a4fb, 32'h42270d05, 32'h428a2b4c};
test_label[1118] = '{32'hc1b7d1b7};
test_output[1118] = '{32'h42f29968};
/*############ DEBUG ############
test_input[8944:8951] = '{-40.0277310082, -98.3504524205, -22.9774007329, -26.2546225837, -39.6374015706, 98.3222238176, 41.7627155825, 69.0845651775};
test_label[1118] = '{-22.9774007329};
test_output[1118] = '{121.29962455};
############ END DEBUG ############*/
test_input[8952:8959] = '{32'hc1b4fc58, 32'h428b5f8c, 32'h41894827, 32'hc1695f9a, 32'hc12258bc, 32'h42c25dc6, 32'h4196adc5, 32'hc2a3846d};
test_label[1119] = '{32'hc2a3846d};
test_output[1119] = '{32'h4332f119};
/*############ DEBUG ############
test_input[8952:8959] = '{-22.6232139733, 69.6866172432, 17.1602302688, -14.5858406636, -10.1466637731, 97.1831527713, 18.8348489723, -81.7586414806};
test_label[1119] = '{-81.7586414806};
test_output[1119] = '{178.941794252};
############ END DEBUG ############*/
test_input[8960:8967] = '{32'hc0fd4ca2, 32'hc0494979, 32'h417a9117, 32'h41a8cca8, 32'hc2b85adb, 32'h424c5cab, 32'h42884eeb, 32'h4208e990};
test_label[1120] = '{32'h417a9117};
test_output[1120] = '{32'h4251f990};
/*############ DEBUG ############
test_input[8960:8967] = '{-7.91560477275, -3.14510940866, 15.6604225524, 21.0999302243, -92.1774509441, 51.0904959232, 68.1541351482, 34.2280877492};
test_label[1120] = '{15.6604225524};
test_output[1120] = '{52.4937126346};
############ END DEBUG ############*/
test_input[8968:8975] = '{32'hc2b6fc41, 32'h42a7461f, 32'h4110845e, 32'h42aa14b7, 32'h419f0ff6, 32'hc223bea9, 32'hc273c077, 32'hc2a67a2c};
test_label[1121] = '{32'hc223bea9};
test_output[1121] = '{32'h42fc648c};
/*############ DEBUG ############
test_input[8968:8975] = '{-91.4926806213, 83.6369565496, 9.03231649523, 85.0404607363, 19.8827936964, -40.936191913, -60.9379550226, -83.2386141558};
test_label[1121] = '{-40.936191913};
test_output[1121] = '{126.196377848};
############ END DEBUG ############*/
test_input[8976:8983] = '{32'hc2738a1b, 32'hc2a0c3ec, 32'h41bff0aa, 32'h429ea5c0, 32'h41cb2a78, 32'h420d96c7, 32'hc2aba0c2, 32'hc19d58a1};
test_label[1122] = '{32'h420d96c7};
test_output[1122] = '{32'h422fb4b9};
/*############ DEBUG ############
test_input[8976:8983] = '{-60.8848688715, -80.3826625841, 23.9925117022, 79.3237327699, 25.3957363516, 35.397244979, -85.8139764524, -19.6682766775};
test_label[1122] = '{35.397244979};
test_output[1122] = '{43.926487791};
############ END DEBUG ############*/
test_input[8984:8991] = '{32'hc1ee483f, 32'hc26a160c, 32'h424a10ca, 32'h41f23032, 32'hc03f7d0c, 32'hc2bee921, 32'h42b06952, 32'hc25fb604};
test_label[1123] = '{32'h424a10ca};
test_output[1123] = '{32'h4216c1da};
/*############ DEBUG ############
test_input[8984:8991] = '{-29.7852770458, -58.521530504, 50.5163963716, 30.2735328361, -2.99200721743, -95.4553289328, 88.2057044823, -55.9277498944};
test_label[1123] = '{50.5163963716};
test_output[1123] = '{37.6893081107};
############ END DEBUG ############*/
test_input[8992:8999] = '{32'hc23e6194, 32'h4159d189, 32'h420bcfd2, 32'hc18d7cae, 32'hc298c662, 32'hc26fc361, 32'hc281cae8, 32'hc174c897};
test_label[1124] = '{32'h4159d189};
test_output[1124] = '{32'h41aab6df};
/*############ DEBUG ############
test_input[8992:8999] = '{-47.5952920507, 13.613656347, 34.9529483017, -17.6858782135, -76.3874648974, -59.9407988518, -64.8963029571, -15.2989717503};
test_label[1124] = '{13.613656347};
test_output[1124] = '{21.3392919552};
############ END DEBUG ############*/
test_input[9000:9007] = '{32'h427a90a3, 32'h4182e04b, 32'h417a6dae, 32'h421bd57d, 32'hc2757573, 32'h4180c0a3, 32'hc1930cdc, 32'hc26fa2d4};
test_label[1125] = '{32'hc2757573};
test_output[1125] = '{32'h42f8030b};
/*############ DEBUG ############
test_input[9000:9007] = '{62.6412453386, 16.3595182331, 15.6517769761, 38.9584845221, -61.364694907, 16.0940609475, -18.3812786304, -59.9090107892};
test_label[1125] = '{-61.364694907};
test_output[1125] = '{124.005940246};
############ END DEBUG ############*/
test_input[9008:9015] = '{32'h4292172c, 32'h41e08db8, 32'hc202e5c8, 32'hbe390474, 32'h426cae48, 32'h41e62245, 32'h427d106c, 32'hc21888b2};
test_label[1126] = '{32'h41e62245};
test_output[1126] = '{32'h42311d44};
/*############ DEBUG ############
test_input[9008:9015] = '{73.0452550737, 28.0691991766, -32.7243955784, -0.180681045883, 59.1701973447, 28.7667336756, 63.2660352906, -38.1334932728};
test_label[1126] = '{28.7667336756};
test_output[1126] = '{44.2785789546};
############ END DEBUG ############*/
test_input[9016:9023] = '{32'h42adecb1, 32'hc2210a1c, 32'hc2841000, 32'hc1f2a06d, 32'hc2725a1c, 32'hc293bf04, 32'h4211de00, 32'hc148eb9e};
test_label[1127] = '{32'h4211de00};
test_output[1127] = '{32'h4249fb63};
/*############ DEBUG ############
test_input[9016:9023] = '{86.9622883995, -40.2598715113, -66.0312496934, -30.3283328779, -60.5879969215, -73.8730752675, 36.4667951521, -12.5575233376};
test_label[1127] = '{36.4667951521};
test_output[1127] = '{50.4954932474};
############ END DEBUG ############*/
test_input[9024:9031] = '{32'h412de708, 32'hc226d33e, 32'hc2aaa9b6, 32'hc2b15dfc, 32'hc16c70a0, 32'h4245ad56, 32'h427f73d0, 32'hc19bf48d};
test_label[1128] = '{32'hc19bf48d};
test_output[1128] = '{32'h42a6b70b};
/*############ DEBUG ############
test_input[9024:9031] = '{10.8689037658, -41.7062909271, -85.3314676324, -88.6835605253, -14.777496567, 49.4192736231, 63.8630983349, -19.4944098792};
test_label[1128] = '{-19.4944098792};
test_output[1128] = '{83.3575087476};
############ END DEBUG ############*/
test_input[9032:9039] = '{32'h429d386e, 32'h42651ce1, 32'hc1538ece, 32'hc12c9c38, 32'hc2b04651, 32'hc1f71757, 32'hc1e15695, 32'hc2a9fbb8};
test_label[1129] = '{32'h429d386e};
test_output[1129] = '{32'h30158b10};
/*############ DEBUG ############
test_input[9032:9039] = '{78.6102110257, 57.2782037259, -13.2223641324, -10.7881396024, -88.1373360811, -30.8863964397, -28.1672765125, -84.9916373531};
test_label[1129] = '{78.6102110257};
test_output[1129] = '{5.44035039388e-10};
############ END DEBUG ############*/
test_input[9040:9047] = '{32'hc20206da, 32'h3fab47c8, 32'hc23a271b, 32'hc1172063, 32'h42a2bec7, 32'h41c733b5, 32'h410b263f, 32'h408f235b};
test_label[1130] = '{32'h410b263f};
test_output[1130] = '{32'h429159ff};
/*############ DEBUG ############
test_input[9040:9047] = '{-32.5066896327, 1.3381280774, -46.5381884383, -9.44540738505, 81.3726096763, 24.9002467446, 8.69683785591, 4.47306601585};
test_label[1130] = '{8.69683785591};
test_output[1130] = '{72.6757718204};
############ END DEBUG ############*/
test_input[9048:9055] = '{32'hc1b4d6aa, 32'h423913cf, 32'h421963bc, 32'hc2acf10f, 32'h40e1227d, 32'hc1bfdf60, 32'h428f0d14, 32'hbf13786e};
test_label[1131] = '{32'hc2acf10f};
test_output[1131] = '{32'h431dff12};
/*############ DEBUG ############
test_input[9048:9055] = '{-22.6048164596, 46.2693433505, 38.3473973387, -86.4708181614, 7.03546010915, -23.9840699855, 71.5255452859, -0.576056353004};
test_label[1131] = '{-86.4708181614};
test_output[1131] = '{157.996363447};
############ END DEBUG ############*/
test_input[9056:9063] = '{32'hc0e74f45, 32'h42a0f868, 32'h4193bde8, 32'hc20c408c, 32'hc232d835, 32'hc29333cf, 32'h41e71596, 32'hc21d64c9};
test_label[1132] = '{32'h42a0f868};
test_output[1132] = '{32'h80000000};
/*############ DEBUG ############
test_input[9056:9063] = '{-7.22842663717, 80.4851665474, 18.4677285463, -35.063034316, -44.7111400727, -73.6011891739, 28.8855397246, -39.3484247209};
test_label[1132] = '{80.4851665474};
test_output[1132] = '{-0.0};
############ END DEBUG ############*/
test_input[9064:9071] = '{32'h4182c7f7, 32'h428ec826, 32'hc2327d20, 32'hc2c2ef23, 32'h41afbc43, 32'h421d6031, 32'h40e35bce, 32'h42acd3c4};
test_label[1133] = '{32'h421d6031};
test_output[1133] = '{32'h423c4758};
/*############ DEBUG ############
test_input[9064:9071] = '{16.3476384404, 71.3909123436, -44.6221914713, -97.4670658592, 21.966924677, 39.343937222, 7.10495666592, 86.4136075473};
test_label[1133] = '{39.343937222};
test_output[1133] = '{47.0696706243};
############ END DEBUG ############*/
test_input[9072:9079] = '{32'h42b5957f, 32'hc1542d61, 32'h420679ad, 32'hc11913df, 32'h42961841, 32'hc2191531, 32'hc27d7d35, 32'hc2ac112c};
test_label[1134] = '{32'h420679ad};
test_output[1134] = '{32'h4264b152};
/*############ DEBUG ############
test_input[9072:9079] = '{90.7919871561, -13.2610785431, 33.6188228342, -9.5673510216, 75.0473729075, -38.2706959246, -63.3722722216, -86.0335352444};
test_label[1134] = '{33.6188228342};
test_output[1134] = '{57.1731644672};
############ END DEBUG ############*/
test_input[9080:9087] = '{32'hc21eba96, 32'hc1facaff, 32'h41c2b3f5, 32'h42a9117b, 32'h42392c1e, 32'hc19a8010, 32'h411dc138, 32'hc269eb89};
test_label[1135] = '{32'hc19a8010};
test_output[1135] = '{32'h42cfb17f};
/*############ DEBUG ############
test_input[9080:9087] = '{-39.682212327, -31.3491189608, 24.3378703567, 84.534144347, 46.2930850541, -19.3125313535, 9.85967216044, -58.4800129332};
test_label[1135] = '{-19.3125313535};
test_output[1135] = '{103.846675701};
############ END DEBUG ############*/
test_input[9088:9095] = '{32'hc20d911d, 32'h42afecd9, 32'h4221ae39, 32'h40c3324a, 32'h42697bd2, 32'hc2749954, 32'hc0671b59, 32'h421b1835};
test_label[1136] = '{32'h40c3324a};
test_output[1136] = '{32'h42a3b9b4};
/*############ DEBUG ############
test_input[9088:9095] = '{-35.391711191, 87.9625904378, 40.4201404438, 6.09988862165, 58.3709176552, -61.1497327896, -3.61104407221, 38.7736412239};
test_label[1136] = '{6.09988862165};
test_output[1136] = '{81.8627018161};
############ END DEBUG ############*/
test_input[9096:9103] = '{32'h428951aa, 32'h42a146f6, 32'hc2446151, 32'hc1345a89, 32'h41821460, 32'h4144ccd0, 32'h4207d63a, 32'hc2c0832d};
test_label[1137] = '{32'hc1345a89};
test_output[1137] = '{32'h42b7d248};
/*############ DEBUG ############
test_input[9096:9103] = '{68.6595027478, 80.6385922863, -49.0950357534, -11.2721034936, 16.2599493083, 12.3000032062, 33.9592058406, -96.256206357};
test_label[1137] = '{-11.2721034936};
test_output[1137] = '{91.9107020539};
############ END DEBUG ############*/
test_input[9104:9111] = '{32'h429639e4, 32'hc2b2af9a, 32'hc1b0925d, 32'hc20e6b9f, 32'hc2197705, 32'h41bd7a28, 32'h428ba743, 32'h41838440};
test_label[1138] = '{32'hc1b0925d};
test_output[1138] = '{32'h42c26111};
/*############ DEBUG ############
test_input[9104:9111] = '{75.1130677964, -89.3429715014, -22.0714672894, -35.605100205, -38.3662293215, 23.6846471407, 69.8266803022, 16.4395756055};
test_label[1138] = '{-22.0714672894};
test_output[1138] = '{97.1895823336};
############ END DEBUG ############*/
test_input[9112:9119] = '{32'hc23fe384, 32'hc294c508, 32'h41fecfb0, 32'hc2a1ec48, 32'hc23bdec2, 32'h42b5d51a, 32'h4297850a, 32'h42786cd1};
test_label[1139] = '{32'hc294c508};
test_output[1139] = '{32'h43254d11};
/*############ DEBUG ############
test_input[9112:9119] = '{-47.9721827351, -74.3848255413, 31.8514097771, -80.961489098, -46.9675383004, 90.916215578, 75.7598405928, 62.106265065};
test_label[1139] = '{-74.3848255413};
test_output[1139] = '{165.301041381};
############ END DEBUG ############*/
test_input[9120:9127] = '{32'hc0f00b1a, 32'h426ac507, 32'hc1aa6e69, 32'hc0a5033c, 32'h42971b5a, 32'h42528d7a, 32'hc28afb60, 32'hc1a0babf};
test_label[1140] = '{32'hc1aa6e69};
test_output[1140] = '{32'h42c1b6f4};
/*############ DEBUG ############
test_input[9120:9127] = '{-7.5013551252, 58.6924090404, -21.3039120691, -5.15664475736, 75.5534218789, 52.6381593654, -69.4909680695, -20.0911853597};
test_label[1140] = '{-21.3039120691};
test_output[1140] = '{96.8573339957};
############ END DEBUG ############*/
test_input[9128:9135] = '{32'hc2c145af, 32'h41c93163, 32'hc2b04f7b, 32'h422e29d8, 32'h42044ff8, 32'hc2641193, 32'h40a7cd81, 32'h428b21b9};
test_label[1141] = '{32'hc2c145af};
test_output[1141] = '{32'h432633b4};
/*############ DEBUG ############
test_input[9128:9135] = '{-96.6360998738, 25.1491149032, -88.1552374712, 43.5408641187, 33.0780946657, -57.0171637491, 5.24383599545, 69.5658654872};
test_label[1141] = '{-96.6360998738};
test_output[1141] = '{166.201965361};
############ END DEBUG ############*/
test_input[9136:9143] = '{32'hc2ad3215, 32'h40c8cd2d, 32'h4259ee70, 32'h4287cfc5, 32'h4273a3d2, 32'hc21702d8, 32'h42486430, 32'h428931bd};
test_label[1142] = '{32'hc2ad3215};
test_output[1142] = '{32'h431b99f1};
/*############ DEBUG ############
test_input[9136:9143] = '{-86.5978134379, 6.27504575209, 54.482850955, 67.9057969955, 60.909981566, -37.7527762442, 50.0978405819, 68.5971480194};
test_label[1142] = '{-86.5978134379};
test_output[1142] = '{155.601331697};
############ END DEBUG ############*/
test_input[9144:9151] = '{32'h4296f5b0, 32'hc281a841, 32'h412ee89b, 32'h4264641b, 32'hc2af9bf6, 32'h429a2783, 32'hc2473e7a, 32'h42b85f72};
test_label[1143] = '{32'hc2af9bf6};
test_output[1143] = '{32'h4333fdb4};
/*############ DEBUG ############
test_input[9144:9151] = '{75.4798573884, -64.8286222444, 10.9317882878, 57.0977609733, -87.8046079275, 77.0771684903, -49.811012714, 92.1864142174};
test_label[1143] = '{-87.8046079275};
test_output[1143] = '{179.991022475};
############ END DEBUG ############*/
test_input[9152:9159] = '{32'h4228ffcb, 32'h41f997ab, 32'h42521fd8, 32'h42addc06, 32'h42934d2c, 32'h41d40e9b, 32'hc249f8ba, 32'hc29f6e55};
test_label[1144] = '{32'hc29f6e55};
test_output[1144] = '{32'h4326a52e};
/*############ DEBUG ############
test_input[9152:9159] = '{42.2497962781, 31.1990559329, 52.5310964467, 86.9297358956, 73.6507242965, 26.5071315718, -50.49289842, -79.7154922076};
test_label[1144] = '{-79.7154922076};
test_output[1144] = '{166.645229813};
############ END DEBUG ############*/
test_input[9160:9167] = '{32'hc2ba6380, 32'hc1123480, 32'h428ba81e, 32'hc2bcba49, 32'h402d0e4c, 32'h42aacd9f, 32'h42263bfe, 32'h429e8d29};
test_label[1145] = '{32'h402d0e4c};
test_output[1145] = '{32'h42a5664b};
/*############ DEBUG ############
test_input[9160:9167] = '{-93.1943372756, -9.13781732333, 69.8283506774, -94.3638344113, 2.70399770135, 85.4016066649, 41.5585860523, 79.2757050952};
test_label[1145] = '{2.70399770135};
test_output[1145] = '{82.6997922707};
############ END DEBUG ############*/
test_input[9168:9175] = '{32'h41eacd5a, 32'h4229d965, 32'hc264e8e0, 32'h42bd44c1, 32'hc23cd5ab, 32'hc2858023, 32'h41d4a7c3, 32'hc2863b0d};
test_label[1146] = '{32'hc2858023};
test_output[1146] = '{32'h43216272};
/*############ DEBUG ############
test_input[9168:9175] = '{29.3502686484, 42.4622975659, -57.2274176764, 94.6342859989, -47.2086597532, -66.750265025, 26.5819139679, -67.1153360009};
test_label[1146] = '{-66.750265025};
test_output[1146] = '{161.384551024};
############ END DEBUG ############*/
test_input[9176:9183] = '{32'h42c38edf, 32'h4152b35b, 32'hc25d3cc4, 32'h4289a858, 32'hc2475283, 32'h425508c9, 32'h42bc8fcf, 32'hc2a712d4};
test_label[1147] = '{32'h42c38edf};
test_output[1147] = '{32'h3cf427bd};
/*############ DEBUG ############
test_input[9176:9183] = '{97.7790486578, 13.1687876498, -55.3093418723, 68.8287938189, -49.830577435, 53.2585789709, 94.2808785563, -83.5367761659};
test_label[1147] = '{97.7790486578};
test_output[1147] = '{0.0298041043473};
############ END DEBUG ############*/
test_input[9184:9191] = '{32'h42b027b5, 32'h40a94b27, 32'hc1f58239, 32'hc1daf105, 32'hc2c7fdb2, 32'h42059350, 32'h42b1b200, 32'h4246d774};
test_label[1148] = '{32'h40a94b27};
test_output[1148] = '{32'h42a7e01a};
/*############ DEBUG ############
test_input[9184:9191] = '{88.0775513554, 5.29042382299, -30.6885844665, -27.3676847436, -99.9954953478, 33.3938586012, 88.8476583136, 49.7104017438};
test_label[1148] = '{5.29042382299};
test_output[1148] = '{83.9376986963};
############ END DEBUG ############*/
test_input[9192:9199] = '{32'h42c65a0f, 32'h425771b9, 32'h4130dd3a, 32'h42a2355f, 32'h417ac5ea, 32'hc29f183a, 32'h42b16c5c, 32'hc25e3f6e};
test_label[1149] = '{32'h425771b9};
test_output[1149] = '{32'h4235426c};
/*############ DEBUG ############
test_input[9192:9199] = '{99.1758952889, 53.8610572254, 11.0540103319, 81.1042425963, 15.6733188922, -79.5473211753, 88.7116410031, -55.5619435666};
test_label[1149] = '{53.8610572254};
test_output[1149] = '{45.3148666159};
############ END DEBUG ############*/
test_input[9200:9207] = '{32'h42ba5cba, 32'h42b12d1d, 32'hc27e23a3, 32'hc28bc98e, 32'hc1e9bd0b, 32'h414206b5, 32'h42ad08fb, 32'h40e8431b};
test_label[1150] = '{32'hc28bc98e};
test_output[1150] = '{32'h4323160a};
/*############ DEBUG ############
test_input[9200:9207] = '{93.1811039904, 88.588109879, -63.5348004152, -69.8936581801, -29.2173066524, 12.126637206, 86.5175423674, 7.25819162897};
test_label[1150] = '{-69.8936581801};
test_output[1150] = '{163.086096787};
############ END DEBUG ############*/
test_input[9208:9215] = '{32'h427f3144, 32'h41849fd8, 32'h42241866, 32'h418395c4, 32'h4259f068, 32'hc29594c5, 32'h42266709, 32'hc24db383};
test_label[1151] = '{32'h4259f068};
test_output[1151] = '{32'h411503ce};
/*############ DEBUG ############
test_input[9208:9215] = '{63.7981105414, 16.5780491626, 41.0238282964, 16.4481286408, 54.4847714517, -74.790569158, 41.6006197564, -51.4253030681};
test_label[1151] = '{54.4847714517};
test_output[1151] = '{9.31342929885};
############ END DEBUG ############*/
test_input[9216:9223] = '{32'hc198f0dd, 32'h4298633b, 32'h404a9a59, 32'hc1e8ec06, 32'h4241beab, 32'hc196b8b2, 32'hc29b2336, 32'hc1275250};
test_label[1152] = '{32'hc1e8ec06};
test_output[1152] = '{32'h42d29e3c};
/*############ DEBUG ############
test_input[9216:9223] = '{-19.1176086181, 76.1938072044, 3.16567052257, -29.1152452522, 48.4362003031, -18.8401826895, -77.5687708893, -10.4575962362};
test_label[1152] = '{-29.1152452522};
test_output[1152] = '{105.309052457};
############ END DEBUG ############*/
test_input[9224:9231] = '{32'h428d7d37, 32'h420a6c87, 32'h42c06cf5, 32'hc28c5a9f, 32'h4256fdda, 32'h429522f9, 32'h410c29e5, 32'h42b5ba57};
test_label[1153] = '{32'h410c29e5};
test_output[1153] = '{32'h42aeea26};
/*############ DEBUG ############
test_input[9224:9231] = '{70.7445568792, 34.6059826512, 96.2128094725, -70.1769926372, 53.7479002433, 74.5683079216, 8.76022794404, 90.8639463735};
test_label[1153] = '{8.76022794404};
test_output[1153] = '{87.4573238187};
############ END DEBUG ############*/
test_input[9232:9239] = '{32'h422b8a12, 32'hc28c559a, 32'hc25f7fa1, 32'hc2b09f23, 32'hc23b6c9d, 32'hc24e55cf, 32'hc0b0ad9f, 32'hc2a91823};
test_label[1154] = '{32'hc24e55cf};
test_output[1154] = '{32'h42bceff1};
/*############ DEBUG ############
test_input[9232:9239] = '{42.8848356046, -70.1671882785, -55.8746365466, -88.310811663, -46.8560658198, -51.583796171, -5.52119410031, -84.5471454768};
test_label[1154] = '{-51.583796171};
test_output[1154] = '{94.4686317756};
############ END DEBUG ############*/
test_input[9240:9247] = '{32'h4198a0a0, 32'h42a176b6, 32'h426faa42, 32'hc231d74a, 32'hc19f5e6c, 32'hc277595d, 32'h4297df30, 32'hc0f51588};
test_label[1155] = '{32'hc0f51588};
test_output[1155] = '{32'h42b0cc45};
/*############ DEBUG ############
test_input[9240:9247] = '{19.0784311011, 80.73185598, 59.9162685957, -44.4602417466, -19.9211040778, -61.8372698241, 75.9359163747, -7.65887838245};
test_label[1155] = '{-7.65887838245};
test_output[1155] = '{88.3989636408};
############ END DEBUG ############*/
test_input[9248:9255] = '{32'hc164ff15, 32'hc28c8eb8, 32'hc20c4b3a, 32'hc231d986, 32'hc2945738, 32'hc2b7d2e7, 32'hbeb37826, 32'hc0f4bebf};
test_label[1156] = '{32'hc0f4bebf};
test_output[1156] = '{32'h40e98cca};
/*############ DEBUG ############
test_input[9248:9255] = '{-14.3122763525, -70.2787450521, -35.0734647885, -44.4624245861, -74.1703523042, -91.9119186363, -0.350526032566, -7.64828456745};
test_label[1156] = '{-7.64828456745};
test_output[1156] = '{7.29843622382};
############ END DEBUG ############*/
test_input[9256:9263] = '{32'hbf206c93, 32'h41dc641a, 32'hc28d670c, 32'h42bec56b, 32'hc29f5619, 32'h428b1fa3, 32'h40f7141b, 32'hc29132f8};
test_label[1157] = '{32'h428b1fa3};
test_output[1157] = '{32'h41ce971f};
/*############ DEBUG ############
test_input[9256:9263] = '{-0.626656731486, 27.5488768638, -70.7012625278, 95.3855829941, -79.6681569555, 69.5617930391, 7.72120415617, -72.599550403};
test_label[1157] = '{69.5617930391};
test_output[1157] = '{25.823789955};
############ END DEBUG ############*/
test_input[9264:9271] = '{32'h42b83ab2, 32'h41cdfb0f, 32'hc2a8d3d4, 32'h428d1422, 32'h41037d21, 32'hc11bcdf2, 32'h429cb44d, 32'hc29b244e};
test_label[1158] = '{32'h42b83ab2};
test_output[1158] = '{32'h358d957c};
/*############ DEBUG ############
test_input[9264:9271] = '{92.114637934, 25.7475876759, -84.4137268032, 70.539321392, 8.21804898628, -9.73777922289, 78.3521528474, -77.5709092796};
test_label[1158] = '{92.114637934};
test_output[1158] = '{1.0548824862e-06};
############ END DEBUG ############*/
test_input[9272:9279] = '{32'h40d5adf0, 32'hc2289038, 32'h41c9c985, 32'hc1f06173, 32'h41202494, 32'h41f90b7b, 32'h42487456, 32'hc2a2a33b};
test_label[1159] = '{32'hc2289038};
test_output[1159] = '{32'h42b88247};
/*############ DEBUG ############
test_input[9272:9279] = '{6.67748263963, -42.1408389726, 25.2233987936, -30.0475832642, 10.0089298836, 31.1306058848, 50.1136085992, -81.3188125773};
test_label[1159] = '{-42.1408389726};
test_output[1159] = '{92.2544475775};
############ END DEBUG ############*/
test_input[9280:9287] = '{32'h42888129, 32'hc28a0364, 32'hc161691c, 32'hc2172092, 32'hc188e33e, 32'hc2443566, 32'hc03b807f, 32'hc2497014};
test_label[1160] = '{32'hc2443566};
test_output[1160] = '{32'h42ea9bdc};
/*############ DEBUG ############
test_input[9280:9287] = '{68.2522693258, -69.0066224785, -14.0881613466, -37.7818071333, -17.1109590068, -49.0521469335, -2.92971780579, -50.3594518771};
test_label[1160] = '{-49.0521469335};
test_output[1160] = '{117.304416259};
############ END DEBUG ############*/
test_input[9288:9295] = '{32'h42a470e3, 32'h428a96dd, 32'h42be0177, 32'hc11e26be, 32'h42b42b48, 32'h428e5b17, 32'h41ff6b39, 32'hc25c3924};
test_label[1161] = '{32'h428a96dd};
test_output[1161] = '{32'h41cdb955};
/*############ DEBUG ############
test_input[9288:9295] = '{82.2204808447, 69.2946533129, 95.0028596046, -9.88445887256, 90.0845351145, 71.1779072113, 31.9273551148, -55.0558026361};
test_label[1161] = '{69.2946533129};
test_output[1161] = '{25.7154938536};
############ END DEBUG ############*/
test_input[9296:9303] = '{32'h429a51b6, 32'hc1981c08, 32'hc25a3c4a, 32'hc28ae9fe, 32'h42131e2c, 32'hc26a73a0, 32'h425d78d0, 32'h418deaca};
test_label[1162] = '{32'hc25a3c4a};
test_output[1162] = '{32'h4303b7ee};
/*############ DEBUG ############
test_input[9296:9303] = '{77.1595934077, -19.0136874288, -54.5588760445, -69.4570193467, 36.7794636841, -58.6129151447, 55.3679825478, 17.7396433752};
test_label[1162] = '{-54.5588760445};
test_output[1162] = '{131.718469453};
############ END DEBUG ############*/
test_input[9304:9311] = '{32'hc25f3a6a, 32'hc209c81a, 32'h42742739, 32'hc2b4c38e, 32'h41ed6610, 32'h427d7087, 32'hc1e2a337, 32'hc2243131};
test_label[1163] = '{32'hc1e2a337};
test_output[1163] = '{32'h42b790fd};
/*############ DEBUG ############
test_input[9304:9311] = '{-55.8070466678, -34.4454128536, 61.038302034, -90.3819435269, 29.6748354669, 63.3598910484, -28.3296946564, -41.0480391167};
test_label[1163] = '{-28.3296946564};
test_output[1163] = '{91.7831831018};
############ END DEBUG ############*/
test_input[9312:9319] = '{32'h423d0697, 32'h424b42f7, 32'hc2488c71, 32'hc1594ceb, 32'hc15d530a, 32'h42b8c2d7, 32'hc22f1ddf, 32'hc2c1587f};
test_label[1164] = '{32'hc15d530a};
test_output[1164] = '{32'h42d46d38};
/*############ DEBUG ############
test_input[9312:9319] = '{47.256435252, 50.8153970729, -50.137150146, -13.5812787616, -13.8327732439, 92.380547679, -43.7791720991, -96.6728466547};
test_label[1164] = '{-13.8327732439};
test_output[1164] = '{106.213320923};
############ END DEBUG ############*/
test_input[9320:9327] = '{32'hc2288c1f, 32'hc2690181, 32'h41d6621c, 32'hc293f93e, 32'hc29fce22, 32'hc20fc674, 32'h42968964, 32'hc29775a1};
test_label[1165] = '{32'hc2690181};
test_output[1165] = '{32'h43058512};
/*############ DEBUG ############
test_input[9320:9327] = '{-42.1368355568, -58.2514702275, 26.7979051592, -73.9868019632, -79.9026007816, -35.9438021325, 75.268341593, -75.7297421146};
test_label[1165] = '{-58.2514702275};
test_output[1165] = '{133.519811821};
############ END DEBUG ############*/
test_input[9328:9335] = '{32'h42626176, 32'h4224d72c, 32'h4207c54b, 32'hc2bba8fd, 32'h42247829, 32'h4224461e, 32'h42c034cc, 32'h42b60d69};
test_label[1166] = '{32'h4207c54b};
test_output[1166] = '{32'h4278aaab};
/*############ DEBUG ############
test_input[9328:9335] = '{56.5951785915, 41.210129134, 33.9426698832, -93.8300589738, 41.1173426824, 41.06847296, 96.1031196927, 91.0261933153};
test_label[1166] = '{33.9426698832};
test_output[1166] = '{62.1666694833};
############ END DEBUG ############*/
test_input[9336:9343] = '{32'hc21ea3fe, 32'h41c0f30e, 32'hc0fcbb7f, 32'h404a5f7a, 32'hc2245c2d, 32'hc1c3e3ed, 32'h4211b8e2, 32'h42a29bd5};
test_label[1167] = '{32'h42a29bd5};
test_output[1167] = '{32'h80000000};
/*############ DEBUG ############
test_input[9336:9343] = '{-39.6601468744, 24.1186793897, -7.89788752571, 3.16207742772, -41.0900146234, -24.4862909547, 36.4305478215, 81.3043601194};
test_label[1167] = '{81.3043601194};
test_output[1167] = '{-0.0};
############ END DEBUG ############*/
test_input[9344:9351] = '{32'h424cb8ee, 32'hc1d7f657, 32'hc1dd1855, 32'h422d2750, 32'hc2962bc0, 32'hc2a49160, 32'hc170d9c9, 32'h42575d97};
test_label[1168] = '{32'hc1dd1855};
test_output[1168] = '{32'h42a3177b};
/*############ DEBUG ############
test_input[9344:9351] = '{51.180593611, -26.9952827667, -27.6368807596, 43.2883913025, -75.0854478369, -82.2839350747, -15.0531706698, 53.8413974804};
test_label[1168] = '{-27.6368807596};
test_output[1168] = '{81.5458603715};
############ END DEBUG ############*/
test_input[9352:9359] = '{32'hc14fd424, 32'hc2a55342, 32'hc2bcddbb, 32'h419c2c20, 32'h429b09c1, 32'h4064f351, 32'h4273d9dc, 32'hc24e5da8};
test_label[1169] = '{32'h419c2c20};
test_output[1169] = '{32'h4267fd73};
/*############ DEBUG ############
test_input[9352:9359] = '{-12.9892922171, -82.6626159198, -94.4330646531, 19.5215450905, 77.5190534841, 3.57735085723, 60.9627545489, -51.5914622674};
test_label[1169] = '{19.5215450905};
test_output[1169] = '{57.9975084582};
############ END DEBUG ############*/
test_input[9360:9367] = '{32'hbf1c3d0f, 32'h422bb486, 32'h4170ae1c, 32'h4208fe9a, 32'h4263a54e, 32'h42962270, 32'h41b1dd0d, 32'h42037356};
test_label[1170] = '{32'h4208fe9a};
test_output[1170] = '{32'h42234645};
/*############ DEBUG ############
test_input[9360:9367] = '{-0.610306704853, 42.9262924257, 15.0425073434, 34.2486327181, 56.9114305915, 75.0672571524, 22.2329342623, 32.8626323783};
test_label[1170] = '{34.2486327181};
test_output[1170] = '{40.8186244472};
############ END DEBUG ############*/
test_input[9368:9375] = '{32'hc2b528cc, 32'hc1b125cf, 32'hc29ace21, 32'hc29dbb21, 32'hc26ebb86, 32'h429a8e47, 32'hc26e1442, 32'h4295152a};
test_label[1171] = '{32'hc1b125cf};
test_output[1171] = '{32'h42c6f7e0};
/*############ DEBUG ############
test_input[9368:9375] = '{-90.5796816042, -22.1434609059, -77.4025964801, -78.8654858122, -59.6831292478, 77.2778869812, -59.5197843935, 74.5413336807};
test_label[1171] = '{-22.1434609059};
test_output[1171] = '{99.4841285693};
############ END DEBUG ############*/
test_input[9376:9383] = '{32'h427b6364, 32'hc27fdcd4, 32'h42c05df4, 32'h427b723d, 32'hc2b79c10, 32'h42b4d193, 32'h42bdabba, 32'hc25dbb24};
test_label[1172] = '{32'hc25dbb24};
test_output[1172] = '{32'h4317d981};
/*############ DEBUG ############
test_input[9376:9383] = '{62.8470602415, -63.9656510922, 96.1835012964, 62.8615605307, -91.804809694, 90.4093212731, 94.8354004306, -55.4327541687};
test_label[1172] = '{-55.4327541687};
test_output[1172] = '{151.849618463};
############ END DEBUG ############*/
test_input[9384:9391] = '{32'h422c6b5a, 32'hbef02c17, 32'h42ba60a3, 32'hc29f9522, 32'hc2b8b03f, 32'h41df4ab4, 32'hc2885d1a, 32'hc1e73cad};
test_label[1173] = '{32'h42ba60a3};
test_output[1173] = '{32'h80000000};
/*############ DEBUG ############
test_input[9384:9391] = '{43.1048357056, -0.469086387335, 93.1887400606, -79.7912712397, -92.3442315806, 27.911475329, -68.1818404198, -28.9046274845};
test_label[1173] = '{93.1887400606};
test_output[1173] = '{-0.0};
############ END DEBUG ############*/
test_input[9392:9399] = '{32'hc1bd6f92, 32'hc1336114, 32'h41b5dfa2, 32'h42bf03db, 32'hc253bd70, 32'hc2c5b662, 32'h42a9de4f, 32'hc181ed4f};
test_label[1174] = '{32'hc2c5b662};
test_output[1174] = '{32'h43425d20};
/*############ DEBUG ############
test_input[9392:9399] = '{-23.6794779773, -11.211200608, 22.7341962726, 95.5075292949, -52.934995922, -98.8562133492, 84.9341934019, -16.2408734353};
test_label[1174] = '{-98.8562133492};
test_output[1174] = '{194.363768233};
############ END DEBUG ############*/
test_input[9400:9407] = '{32'h42b1cd97, 32'h42b1f730, 32'h422aa647, 32'h42482b5c, 32'h42937dea, 32'h423f8e26, 32'h42b2dd77, 32'h418d89e3};
test_label[1175] = '{32'h422aa647};
test_output[1175] = '{32'h423e47f9};
/*############ DEBUG ############
test_input[9400:9407] = '{88.9015461495, 88.9827880201, 42.6623795365, 50.0423425132, 73.7459275113, 47.8888154918, 89.4325512505, 17.6923275765};
test_label[1175] = '{42.6623795365};
test_output[1175] = '{47.5702849499};
############ END DEBUG ############*/
test_input[9408:9415] = '{32'hc29bef2f, 32'hc281b4a7, 32'hc28c1cca, 32'h41035002, 32'hc280e5a4, 32'h3f635326, 32'h41885969, 32'h4265e1a0};
test_label[1176] = '{32'hc29bef2f};
test_output[1176] = '{32'h43077000};
/*############ DEBUG ############
test_input[9408:9415] = '{-77.96715719, -64.8528390465, -70.0562297417, 8.20703305361, -64.4485177956, 0.887987476703, 17.0436571249, 57.470337558};
test_label[1176] = '{-77.96715719};
test_output[1176] = '{135.437494748};
############ END DEBUG ############*/
test_input[9416:9423] = '{32'h424b7f89, 32'h4295ad82, 32'hc2919bdb, 32'hc238325d, 32'hc2b5614b, 32'h415277d9, 32'h42c079b7, 32'hc2970712};
test_label[1177] = '{32'hc2919bdb};
test_output[1177] = '{32'h43290ac9};
/*############ DEBUG ############
test_input[9416:9423] = '{50.874547389, 74.8388855653, -72.8044058748, -46.0491810216, -90.6900245374, 13.1542597805, 96.2377220101, -75.5138058523};
test_label[1177] = '{-72.8044058748};
test_output[1177] = '{169.042127885};
############ END DEBUG ############*/
test_input[9424:9431] = '{32'hc298f42d, 32'h4231deb7, 32'hc2c0c310, 32'h424b35e8, 32'h411337e1, 32'hc26299b0, 32'hc2bab8ab, 32'h41fd4a5f};
test_label[1178] = '{32'h411337e1};
test_output[1178] = '{32'h422669c1};
/*############ DEBUG ############
test_input[9424:9431] = '{-76.4769030905, 44.467494716, -96.3809837348, 50.8026442789, 9.20114183584, -56.6500871038, -93.3606785989, 31.6613138471};
test_label[1178] = '{9.20114183584};
test_output[1178] = '{41.6032737588};
############ END DEBUG ############*/
test_input[9432:9439] = '{32'hc2340170, 32'hc25a9138, 32'h424f425d, 32'h41320c18, 32'h41a537d7, 32'h42ac2fae, 32'h40e0422e, 32'h41127100};
test_label[1179] = '{32'hc25a9138};
test_output[1179] = '{32'h430cbc25};
/*############ DEBUG ############
test_input[9432:9439] = '{-45.0014020984, -54.6418155476, 51.8148096554, 11.1279528101, 20.6522651462, 86.0931214467, 7.0080784376, 9.15258780309};
test_label[1179] = '{-54.6418155476};
test_output[1179] = '{140.734936994};
############ END DEBUG ############*/
test_input[9440:9447] = '{32'h4273dbe3, 32'h428e16c0, 32'hc203cb9f, 32'hc2a07684, 32'hc24ced44, 32'hc292ce5f, 32'hc1510dc4, 32'hc2aad865};
test_label[1180] = '{32'hc1510dc4};
test_output[1180] = '{32'h42a8387e};
/*############ DEBUG ############
test_input[9440:9447] = '{60.9647325724, 71.0444357309, -32.948850273, -80.2314778271, -51.2317030728, -73.4030722039, -13.0658604879, -85.4226482417};
test_label[1180] = '{-13.0658604879};
test_output[1180] = '{84.1103381398};
############ END DEBUG ############*/
test_input[9448:9455] = '{32'h42b82671, 32'h4222b959, 32'hc2b8d8e8, 32'hc0864ead, 32'h429542e5, 32'h42ae7112, 32'h42852c5c, 32'h42c6a0e2};
test_label[1181] = '{32'h42ae7112};
test_output[1181] = '{32'h41418176};
/*############ DEBUG ############
test_input[9448:9455] = '{92.0750800715, 40.68100192, -92.4236432778, -4.19710379639, 74.6306534444, 87.2208371169, 66.5866357404, 99.3142208966};
test_label[1181] = '{87.2208371169};
test_output[1181] = '{12.0941070428};
############ END DEBUG ############*/
test_input[9456:9463] = '{32'hc23846e9, 32'hc2015f41, 32'h41fba0d4, 32'h42817668, 32'hc2018b36, 32'hc22bfb91, 32'hc208b5f7, 32'h42894a7b};
test_label[1182] = '{32'h41fba0d4};
test_output[1182] = '{32'h4214d8c9};
/*############ DEBUG ############
test_input[9456:9463] = '{-46.0692482688, -32.3430214328, 31.4535294345, 64.7312617466, -32.3859488786, -42.9956687566, -34.1777006513, 68.6454732313};
test_label[1182] = '{31.4535294345};
test_output[1182] = '{37.2117035587};
############ END DEBUG ############*/
test_input[9464:9471] = '{32'h409b45e6, 32'h420fd19e, 32'h42a68b43, 32'hc116dde7, 32'hc2bb7437, 32'h4288ad76, 32'hc2aed589, 32'hc297cf63};
test_label[1183] = '{32'h420fd19e};
test_output[1183] = '{32'h423d44e9};
/*############ DEBUG ############
test_input[9464:9471] = '{4.8522823567, 35.9547034459, 83.2719982079, -9.42917549516, -93.726985591, 68.3387871789, -87.4170638426, -75.9050549357};
test_label[1183] = '{35.9547034459};
test_output[1183] = '{47.3172950891};
############ END DEBUG ############*/
test_input[9472:9479] = '{32'hc22f820d, 32'h4240ccc4, 32'hc2647cab, 32'hc2281641, 32'h41a94195, 32'hc2c38468, 32'h405bf466, 32'h415b473b};
test_label[1184] = '{32'h415b473b};
test_output[1184] = '{32'h4209faf6};
/*############ DEBUG ############
test_input[9472:9479] = '{-43.8770039543, 48.1999674925, -57.1217455118, -42.0217340927, 21.1570232245, -97.7586082864, 3.43679177867, 13.7048901688};
test_label[1184] = '{13.7048901688};
test_output[1184] = '{34.4950773238};
############ END DEBUG ############*/
test_input[9480:9487] = '{32'hc031158a, 32'hc22a517f, 32'h4285c024, 32'hc1fc5195, 32'h42addb5f, 32'h4213f32b, 32'hc2c63317, 32'hc0e1b75d};
test_label[1185] = '{32'hc0e1b75d};
test_output[1185] = '{32'h42bbf6d5};
/*############ DEBUG ############
test_input[9480:9487] = '{-2.76693952681, -42.5795864302, 66.8752713076, -31.5398342172, 86.928459616, 36.9874693738, -99.0997863499, -7.05363326581};
test_label[1185] = '{-7.05363326581};
test_output[1185] = '{93.9820928838};
############ END DEBUG ############*/
test_input[9488:9495] = '{32'hc26f4e01, 32'hbfd229e7, 32'hc08b5e86, 32'hc26ecd83, 32'hc2946e74, 32'h41cb185e, 32'hc24dc6cc, 32'h42621c9f};
test_label[1186] = '{32'hc26ecd83};
test_output[1186] = '{32'h42e87511};
/*############ DEBUG ############
test_input[9488:9495] = '{-59.8261768892, -1.64190377663, -4.35528865373, -59.7006937628, -74.2157280102, 25.3868971117, -51.4441386345, 56.5279518798};
test_label[1186] = '{-59.7006937628};
test_output[1186] = '{116.228645643};
############ END DEBUG ############*/
test_input[9496:9503] = '{32'hc27435cf, 32'h41d28be5, 32'hc2937ba4, 32'hc243bb85, 32'h4285b76c, 32'hc1b170dd, 32'h423f2088, 32'h41eb8082};
test_label[1187] = '{32'h4285b76c};
test_output[1187] = '{32'h31b25676};
/*############ DEBUG ############
test_input[9496:9503] = '{-61.0525479918, 26.31830707, -73.7414884358, -48.9331229835, 66.8582424649, -22.1801086667, 47.7817703083, 29.437748072};
test_label[1187] = '{66.8582424649};
test_output[1187] = '{5.19031130534e-09};
############ END DEBUG ############*/
test_input[9504:9511] = '{32'h40a065e8, 32'h420e2599, 32'h42aa4617, 32'h429de2db, 32'hc28e059c, 32'h42b6cdd9, 32'h42264177, 32'hc24c1877};
test_label[1188] = '{32'hc28e059c};
test_output[1188] = '{32'h43226a37};
/*############ DEBUG ############
test_input[9504:9511] = '{5.01243984372, 35.5367154814, 85.1368951389, 78.9430779704, -71.0109589319, 91.4020466313, 41.5639317406, -51.0238897244};
test_label[1188] = '{-71.0109589319};
test_output[1188] = '{162.414909058};
############ END DEBUG ############*/
test_input[9512:9519] = '{32'h42b508a9, 32'h406a984c, 32'hc2ae5e55, 32'h41a6406b, 32'hc2b6abba, 32'hc283054f, 32'hc12a45b5, 32'hc01cdc08};
test_label[1189] = '{32'hc283054f};
test_output[1189] = '{32'h431c06fc};
/*############ DEBUG ############
test_input[9512:9519] = '{90.5169117097, 3.66554543537, -87.1842438054, 20.7814550098, -91.3354070112, -65.5103684023, -10.6420181227, -2.4509297086};
test_label[1189] = '{-65.5103684023};
test_output[1189] = '{156.027280112};
############ END DEBUG ############*/
test_input[9520:9527] = '{32'hc2a94c66, 32'h42985118, 32'h4240f6cb, 32'h426c2f74, 32'h42c5ebfa, 32'h41d650cc, 32'h428836d9, 32'h42073d5c};
test_label[1190] = '{32'h41d650cc};
test_output[1190] = '{32'h429057c7};
/*############ DEBUG ############
test_input[9520:9527] = '{-84.6492169436, 76.1583862187, 48.2410103565, 59.0463413108, 98.9608952155, 26.7894518801, 68.1071230633, 33.8099197775};
test_label[1190] = '{26.7894518801};
test_output[1190] = '{72.1714433356};
############ END DEBUG ############*/
test_input[9528:9535] = '{32'hc24bf4d7, 32'h40c6ac24, 32'h4181223c, 32'hc10d55f7, 32'h42ac0929, 32'hc212fb59, 32'h42b63ac8, 32'hc2348e9e};
test_label[1191] = '{32'h42ac0929};
test_output[1191] = '{32'h40a34be4};
/*############ DEBUG ############
test_input[9528:9535] = '{-50.9891000528, 6.20851335648, 16.1417164734, -8.83348734992, 86.017890367, -36.7454565921, 91.1148075523, -45.1392747846};
test_label[1191] = '{86.017890367};
test_output[1191] = '{5.10301413183};
############ END DEBUG ############*/
test_input[9536:9543] = '{32'h4219abf7, 32'h4182c7d1, 32'hc21830fa, 32'h426f5928, 32'hc2b6479e, 32'hc23fa92d, 32'hc25ebdc7, 32'h425ecfd3};
test_label[1192] = '{32'hc2b6479e};
test_output[1192] = '{32'h4316fe2a};
/*############ DEBUG ############
test_input[9536:9543] = '{38.4179342887, 16.3475674141, -38.0478305473, 59.8370659093, -91.1398737661, -47.9152093177, -55.6853292822, 55.7029536572};
test_label[1192] = '{-91.1398737661};
test_output[1192] = '{150.992829637};
############ END DEBUG ############*/
test_input[9544:9551] = '{32'hc2412ee4, 32'hc2a0a35e, 32'h42622b93, 32'h421ecb17, 32'hc2804a04, 32'hc21b41c3, 32'hc2a5b7d0, 32'hc10f93ac};
test_label[1193] = '{32'hc2a0a35e};
test_output[1193] = '{32'h4308dc94};
/*############ DEBUG ############
test_input[9544:9551] = '{-48.2957919114, -80.3190767556, 56.5425523467, 39.6983284667, -64.1445651886, -38.8142188288, -82.8590097202, -8.97355296062};
test_label[1193] = '{-80.3190767556};
test_output[1193] = '{136.861629151};
############ END DEBUG ############*/
test_input[9552:9559] = '{32'hc220f47a, 32'hc20f17b3, 32'hbf129532, 32'hc2a6499c, 32'h42160d21, 32'h4219d66d, 32'hc2c77166, 32'h41903924};
test_label[1194] = '{32'hc2c77166};
test_output[1194] = '{32'h430a8240};
/*############ DEBUG ############
test_input[9552:9559] = '{-40.2387464493, -35.7731442807, -0.572589038901, -83.1437658078, 37.51282207, 38.4594002943, -99.7214782978, 18.0279001328};
test_label[1194] = '{-99.7214782978};
test_output[1194] = '{138.508790459};
############ END DEBUG ############*/
test_input[9560:9567] = '{32'h41ee7c02, 32'h418caebf, 32'hc27412a0, 32'h42669ef1, 32'hc217f1b9, 32'h429681e7, 32'h42b7e5b2, 32'hc20e0684};
test_label[1195] = '{32'h42669ef1};
test_output[1195] = '{32'h42092c72};
/*############ DEBUG ############
test_input[9560:9567] = '{29.8105507405, 17.5853247534, -61.0181887035, 57.6552166543, -37.9860583379, 75.2537149686, 91.9486206525, -35.5063622945};
test_label[1195] = '{57.6552166543};
test_output[1195] = '{34.2934040544};
############ END DEBUG ############*/
test_input[9568:9575] = '{32'hc0a5b599, 32'hc2038c6b, 32'h41cf4027, 32'hc1b8c149, 32'hc1b0c18b, 32'hc23598d5, 32'h42c00399, 32'h426f5479};
test_label[1196] = '{32'hc23598d5};
test_output[1196] = '{32'h430d6802};
/*############ DEBUG ############
test_input[9568:9575] = '{-5.17841754904, -32.8871251911, 25.906324396, -23.0943771335, -22.0945030591, -45.399251172, 96.007026912, 59.8324944673};
test_label[1196] = '{-45.399251172};
test_output[1196] = '{141.406278084};
############ END DEBUG ############*/
test_input[9576:9583] = '{32'h41ba00af, 32'hc0d96cd4, 32'h42b0ad59, 32'h427c3087, 32'h4275c48a, 32'hc2a56b99, 32'hc246736a, 32'h416dddf9};
test_label[1197] = '{32'h427c3087};
test_output[1197] = '{32'h41ca5458};
/*############ DEBUG ############
test_input[9576:9583] = '{23.2503342475, -6.79453473187, 88.3385727751, 63.0473893378, 61.4419314759, -82.7101510814, -49.6127095089, 14.8666923726};
test_label[1197] = '{63.0473893378};
test_output[1197] = '{25.2911834374};
############ END DEBUG ############*/
test_input[9584:9591] = '{32'hc28f9d4a, 32'hc29df5ab, 32'hc152b8b0, 32'h423f6cd4, 32'h41cd3892, 32'hc2027b3e, 32'hc2c07dea, 32'h4288f6d9};
test_label[1198] = '{32'h41cd3892};
test_output[1198] = '{32'h422b5169};
/*############ DEBUG ############
test_input[9584:9591] = '{-71.8072020153, -78.979823308, -13.1700901623, 47.8562782172, 25.6526230249, -32.6203527709, -96.2459292976, 68.4821259098};
test_label[1198] = '{25.6526230249};
test_output[1198] = '{42.8295028861};
############ END DEBUG ############*/
test_input[9592:9599] = '{32'hc298143c, 32'h40ae7138, 32'h42708be8, 32'hc08d710f, 32'hc2b36159, 32'h407c76f7, 32'h420bcba3, 32'hc1993c67};
test_label[1199] = '{32'hc1993c67};
test_output[1199] = '{32'h429e950e};
/*############ DEBUG ############
test_input[9592:9599] = '{-76.0395231489, 5.45132081549, 60.1366274045, -4.42005097047, -89.6901327284, 3.94476115359, 34.9488622913, -19.1544925445};
test_label[1199] = '{-19.1544925445};
test_output[1199] = '{79.291119949};
############ END DEBUG ############*/
test_input[9600:9607] = '{32'hc2a09309, 32'hc0e10724, 32'hc25b5726, 32'hc249260f, 32'h411a1eb3, 32'hc224242c, 32'hc2a41910, 32'hc2bf87db};
test_label[1200] = '{32'hc25b5726};
test_output[1200] = '{32'h4280ef69};
/*############ DEBUG ############
test_input[9600:9607] = '{-80.2871789836, -7.03212174032, -54.8351059476, -50.2871660809, 9.63249472974, -41.0353236485, -82.0489530756, -95.7653417053};
test_label[1200] = '{-54.8351059476};
test_output[1200] = '{64.4676007353};
############ END DEBUG ############*/
test_input[9608:9615] = '{32'h42bb9ad3, 32'hc1f279f9, 32'hbf0c11d7, 32'hc22ea836, 32'h4280d10a, 32'h412d0714, 32'h42441ec5, 32'h418df946};
test_label[1201] = '{32'hbf0c11d7};
test_output[1201] = '{32'h42bcb2f7};
/*############ DEBUG ############
test_input[9608:9615] = '{93.8023901408, -30.309557289, -0.547147211557, -43.6642689489, 64.4082807482, 10.8142276845, 49.0300471467, 17.7467157333};
test_label[1201] = '{-0.547147211557};
test_output[1201] = '{94.3495373524};
############ END DEBUG ############*/
test_input[9616:9623] = '{32'h4099b861, 32'hc2108b0f, 32'h42bf0ff1, 32'hc23e664f, 32'hc1382be2, 32'h4223d025, 32'h422549fc, 32'hc27b1b3f};
test_label[1202] = '{32'hc23e664f};
test_output[1202] = '{32'h430f218c};
/*############ DEBUG ############
test_input[9616:9623] = '{4.80375728223, -36.1358003961, 95.5311334529, -47.5999109825, -11.5107136664, 40.9532680074, 41.3222516016, -62.7766056182};
test_label[1202] = '{-47.5999109825};
test_output[1202] = '{143.131044435};
############ END DEBUG ############*/
test_input[9624:9631] = '{32'hc2610e1e, 32'h426745aa, 32'hc285efe1, 32'hc2563b4b, 32'hc0877ff5, 32'hbf7d141c, 32'h42c43ecf, 32'h42020ad6};
test_label[1203] = '{32'hbf7d141c};
test_output[1203] = '{32'h42c638f7};
/*############ DEBUG ############
test_input[9624:9631] = '{-56.2637872561, 57.8180294902, -66.9685098395, -53.5579039196, -4.23436970231, -0.988588110322, 98.1226695815, 32.5105805774};
test_label[1203] = '{-0.988588110322};
test_output[1203] = '{99.1112576919};
############ END DEBUG ############*/
test_input[9632:9639] = '{32'h42bf1de2, 32'hc2b4c1fd, 32'hc213ebaf, 32'hc20fba76, 32'h42823d29, 32'hc2022cc6, 32'hc126274c, 32'h420df0cb};
test_label[1204] = '{32'hc20fba76};
test_output[1204] = '{32'h43037d8f};
/*############ DEBUG ############
test_input[9632:9639] = '{95.5583657712, -90.3788814452, -36.9801614472, -35.9320905537, 65.1194530937, -32.5437237942, -10.3845940293, 35.4851485586};
test_label[1204] = '{-35.9320905537};
test_output[1204] = '{131.490456325};
############ END DEBUG ############*/
test_input[9640:9647] = '{32'hc299d7b5, 32'h42a979bd, 32'hc284431b, 32'h4214b51e, 32'h42c05afa, 32'h42bba2a1, 32'h428d4038, 32'h41cdf68c};
test_label[1205] = '{32'hc284431b};
test_output[1205] = '{32'h43226624};
/*############ DEBUG ############
test_input[9640:9647] = '{-76.9213064502, 84.7377725224, -66.1310657683, 37.1768723739, 96.1776921554, 93.8176373855, 70.625429175, 25.7453842635};
test_label[1205] = '{-66.1310657683};
test_output[1205] = '{162.398987774};
############ END DEBUG ############*/
test_input[9648:9655] = '{32'hc215ff9e, 32'h42a3f7f3, 32'h40cafea1, 32'hc291613a, 32'h42173c0b, 32'hc242367e, 32'h429187bc, 32'h42b477e0};
test_label[1206] = '{32'h40cafea1};
test_output[1206] = '{32'h42a7c818};
/*############ DEBUG ############
test_input[9648:9655] = '{-37.4996258877, 81.9842754369, 6.34358268971, -72.6898974208, 37.8086370419, -48.5532167573, 72.7651030283, 90.2341323397};
test_label[1206] = '{6.34358268971};
test_output[1206] = '{83.8908109377};
############ END DEBUG ############*/
test_input[9656:9663] = '{32'h42648b46, 32'h42b61514, 32'hc1214909, 32'hc29159c3, 32'h418079d9, 32'h427646f3, 32'h4188cd7f, 32'hc29866f5};
test_label[1207] = '{32'hc29866f5};
test_output[1207] = '{32'h43273e05};
/*############ DEBUG ############
test_input[9656:9663] = '{57.136007411, 91.0411678274, -10.0803311941, -72.6753124747, 16.0594960681, 61.5692875837, 17.1003406114, -76.2010905631};
test_label[1207] = '{-76.2010905631};
test_output[1207] = '{167.24225839};
############ END DEBUG ############*/
test_input[9664:9671] = '{32'h41550e77, 32'h42be970b, 32'h42bfbe2d, 32'h429074e4, 32'h42976c2c, 32'h42324530, 32'h4270ada1, 32'h42892611};
test_label[1208] = '{32'h41550e77};
test_output[1208] = '{32'h42a600ac};
/*############ DEBUG ############
test_input[9664:9671] = '{13.3160316807, 95.2950093048, 95.8714393171, 72.2282985594, 75.7112763257, 44.567566452, 60.1695612975, 68.5743519236};
test_label[1208] = '{13.3160316807};
test_output[1208] = '{83.0013111588};
############ END DEBUG ############*/
test_input[9672:9679] = '{32'h42ac43bf, 32'hc1dc1cd1, 32'h427e35db, 32'hc29de854, 32'h428e8a80, 32'hc2b7bc88, 32'h4216d705, 32'h4250002b};
test_label[1209] = '{32'hc29de854};
test_output[1209] = '{32'h43251609};
/*############ DEBUG ############
test_input[9672:9679] = '{86.1323128437, -27.5140710134, 63.5525924005, -78.9537677382, 71.2705066164, -91.8682264065, 37.7099813691, 52.0001659235};
test_label[1209] = '{-78.9537677382};
test_output[1209] = '{165.086080933};
############ END DEBUG ############*/
test_input[9680:9687] = '{32'hc205a997, 32'h3f90d882, 32'hc28eab4b, 32'hc20bf58e, 32'h42bb9f9e, 32'h42c72f7e, 32'hc25f31b5, 32'h429cdbfd};
test_label[1210] = '{32'hc20bf58e};
test_output[1210] = '{32'h430695ec};
/*############ DEBUG ############
test_input[9680:9687] = '{-33.4156143801, 1.13160730156, -71.3345584503, -34.98980041, 93.8117530062, 99.5927546924, -55.7985418696, 78.429661704};
test_label[1210] = '{-34.98980041};
test_output[1210] = '{134.585635975};
############ END DEBUG ############*/
test_input[9688:9695] = '{32'h422069e2, 32'hc0a21927, 32'hc283a5ee, 32'hc1981a11, 32'h42989c9e, 32'hc1faf8d7, 32'hc1994a6f, 32'h421d1e5a};
test_label[1211] = '{32'hc1981a11};
test_output[1211] = '{32'h42bea322};
/*############ DEBUG ############
test_input[9688:9695] = '{40.1034002706, -5.06557052838, -65.8240821743, -19.0127286627, 76.3058923727, -31.3715035429, -19.1613447471, 39.2796393809};
test_label[1211] = '{-19.0127286627};
test_output[1211] = '{95.3186210354};
############ END DEBUG ############*/
test_input[9696:9703] = '{32'h4204495b, 32'hc205355e, 32'hc25a601c, 32'hc257e515, 32'h4201e095, 32'hc2acd3e5, 32'hc2a0b4d9, 32'hc1f2aac7};
test_label[1212] = '{32'hc25a601c};
test_output[1212] = '{32'h42b0344f};
/*############ DEBUG ############
test_input[9696:9703] = '{33.0716369877, -33.3021177441, -54.5938582974, -53.9737116036, 32.4693199041, -86.413858867, -80.3532169203, -30.3333864722};
test_label[1212] = '{-54.5938582974};
test_output[1212] = '{88.1021628056};
############ END DEBUG ############*/
test_input[9704:9711] = '{32'h42a7519e, 32'hc2c345cd, 32'h40756254, 32'h3f194bd3, 32'h428eab1a, 32'h42013490, 32'h42b30868, 32'hc23f163b};
test_label[1213] = '{32'h42a7519e};
test_output[1213] = '{32'h40bb8401};
/*############ DEBUG ############
test_input[9704:9711] = '{83.6594121575, -97.6363334354, 3.8341265767, 0.598813215311, 71.3341801861, 32.3013313006, 89.5164202319, -47.7717093801};
test_label[1213] = '{83.6594121575};
test_output[1213] = '{5.85986379274};
############ END DEBUG ############*/
test_input[9712:9719] = '{32'h42acec25, 32'h40bf5f6c, 32'h40fa80bf, 32'h42bdaab0, 32'hc2012534, 32'hc18a098d, 32'h42c1ed85, 32'h41f65fc2};
test_label[1214] = '{32'h40fa80bf};
test_output[1214] = '{32'h42b27ef3};
/*############ DEBUG ############
test_input[9712:9719] = '{86.461218872, 5.9803983863, 7.82821628151, 94.8333707587, -32.286332231, -17.2546633216, 96.9639087106, 30.7967567254};
test_label[1214] = '{7.82821628151};
test_output[1214] = '{89.2479498665};
############ END DEBUG ############*/
test_input[9720:9727] = '{32'h41822d87, 32'h41c57568, 32'hc2776c37, 32'hc2c3aad6, 32'h42ae36c3, 32'h4212e384, 32'hc28800a7, 32'h423f0384};
test_label[1215] = '{32'h41c57568};
test_output[1215] = '{32'h4279b2d2};
/*############ DEBUG ############
test_input[9720:9727] = '{16.2722294549, 24.6823279594, -61.8556804392, -97.8336615538, 87.1069575628, 36.722182249, -68.0012772059, 47.7534325755};
test_label[1215] = '{24.6823279594};
test_output[1215] = '{62.4246296034};
############ END DEBUG ############*/
test_input[9728:9735] = '{32'h425704b0, 32'h4260d4f5, 32'hc2370faf, 32'hc22b7cf4, 32'hc224b1a5, 32'h421cb914, 32'h427a0cd0, 32'hc200a268};
test_label[1216] = '{32'h425704b0};
test_output[1216] = '{32'h410c289f};
/*############ DEBUG ############
test_input[9728:9735] = '{53.7545774789, 56.2079676105, -45.7653154781, -42.8720257701, -41.1734822727, 39.1807392596, 62.5125116995, -32.1586003934};
test_label[1216] = '{53.7545774789};
test_output[1216] = '{8.7599174413};
############ END DEBUG ############*/
test_input[9736:9743] = '{32'hc1ce1e4f, 32'h4282127b, 32'h42955d63, 32'hc2922e4f, 32'hc2c2b700, 32'hc2a9cfbf, 32'h4278d8eb, 32'h4240034e};
test_label[1217] = '{32'h4282127b};
test_output[1217] = '{32'h411a5786};
/*############ DEBUG ############
test_input[9736:9743] = '{-25.7647995253, 65.0360953037, 74.6823950844, -73.0904445753, -97.3574218775, -84.9057513579, 62.2118336249, 48.0032255703};
test_label[1217] = '{65.0360953037};
test_output[1217] = '{9.64636828079};
############ END DEBUG ############*/
test_input[9744:9751] = '{32'hc28e8a76, 32'h422c405b, 32'h42a43290, 32'hc27a454e, 32'hc1ae3100, 32'hc24da205, 32'h4210b3c8, 32'hc2ba0e04};
test_label[1218] = '{32'hc28e8a76};
test_output[1218] = '{32'h43195e83};
/*############ DEBUG ############
test_input[9744:9751] = '{-71.2704301303, 43.0628484237, 82.0987518873, -62.5676812583, -21.7739264162, -51.4082206688, 36.1755674484, -93.0273718318};
test_label[1218] = '{-71.2704301303};
test_output[1218] = '{153.369182018};
############ END DEBUG ############*/
test_input[9752:9759] = '{32'h42c332c6, 32'hc2bb5468, 32'h42097656, 32'h415a37d6, 32'h429d6b96, 32'hc215433c, 32'h425507c0, 32'hc0a171f5};
test_label[1219] = '{32'h415a37d6};
test_output[1219] = '{32'h42a7ebcc};
/*############ DEBUG ############
test_input[9752:9759] = '{97.5991693865, -93.6648581333, 34.365561197, 13.6386321598, 78.7101308488, -37.3156602999, 53.2575698352, -5.04516094391};
test_label[1219] = '{13.6386321598};
test_output[1219] = '{83.9605372331};
############ END DEBUG ############*/
test_input[9760:9767] = '{32'h42a27bc5, 32'hc18001a7, 32'hc298d24c, 32'h4184c54b, 32'hc27761b6, 32'hc2931bbc, 32'hc22bc139, 32'hc2017206};
test_label[1220] = '{32'h42a27bc5};
test_output[1220] = '{32'h80000000};
/*############ DEBUG ############
test_input[9760:9767] = '{81.241737985, -16.0008070475, -76.4107366119, 16.5963350952, -61.8454206302, -73.554169494, -42.9386949293, -32.3613492779};
test_label[1220] = '{81.241737985};
test_output[1220] = '{-0.0};
############ END DEBUG ############*/
test_input[9768:9775] = '{32'h426a71b1, 32'hc217ab0b, 32'hc14a1828, 32'hc2416577, 32'hc180ca9f, 32'h42a92965, 32'h423be5c1, 32'hc27eb982};
test_label[1221] = '{32'hc2416577};
test_output[1221] = '{32'h4304ee10};
/*############ DEBUG ############
test_input[9768:9775] = '{58.6110278586, -37.9170355851, -12.6308978346, -48.3490848717, -16.0989359964, 84.5808450443, 46.9743694373, -63.681161055};
test_label[1221] = '{-48.3490848717};
test_output[1221] = '{132.929929916};
############ END DEBUG ############*/
test_input[9776:9783] = '{32'h425e4a2a, 32'hc28ca730, 32'h41abf285, 32'hc27b8374, 32'h42c26eac, 32'hc21761dc, 32'hc1b46410, 32'h4131cc6f};
test_label[1222] = '{32'hc21761dc};
test_output[1222] = '{32'h43070fcd};
/*############ DEBUG ############
test_input[9776:9783] = '{55.5724268301, -70.3265418239, 21.4934168208, -62.8783738062, 97.2161556294, -37.8455650115, -22.5488579009, 11.1124101193};
test_label[1222] = '{-37.8455650115};
test_output[1222] = '{135.061720641};
############ END DEBUG ############*/
test_input[9784:9791] = '{32'h42107df7, 32'h4281166c, 32'hc2ac76d6, 32'h426de335, 32'hc26800e7, 32'hbf5df4d6, 32'h419a752c, 32'hc291c76f};
test_label[1223] = '{32'h426de335};
test_output[1223] = '{32'h40a28048};
/*############ DEBUG ############
test_input[9784:9791] = '{36.1230107196, 64.5437895572, -86.2321000829, 59.4718813252, -58.0008824776, -0.867017127571, 19.3072120389, -72.8895184374};
test_label[1223] = '{59.4718813252};
test_output[1223] = '{5.07815909779};
############ END DEBUG ############*/
test_input[9792:9799] = '{32'hc0f61b41, 32'hc28dc4cc, 32'hc2943dc1, 32'h42ad3be7, 32'h4286ec53, 32'hc1db7efa, 32'h40bd3f8e, 32'h41df99b4};
test_label[1224] = '{32'hc28dc4cc};
test_output[1224] = '{32'h431d8059};
/*############ DEBUG ############
test_input[9792:9799] = '{-7.69082666128, -70.8843660978, -74.1206135973, 86.6169958114, 67.4615711826, -27.4370000173, 5.91400812287, 27.950049582};
test_label[1224] = '{-70.8843660978};
test_output[1224] = '{157.501361914};
############ END DEBUG ############*/
test_input[9800:9807] = '{32'h41de85fb, 32'h41a95f33, 32'h427c9308, 32'hc2ba7b23, 32'h4291d8bf, 32'h41d402f2, 32'h41ce85ee, 32'hc29b620b};
test_label[1225] = '{32'h41a95f33};
test_output[1225] = '{32'h424f01f3};
/*############ DEBUG ############
test_input[9800:9807] = '{27.8154194564, 21.1714845864, 63.1435835976, -93.2405014254, 72.9233305847, 26.5014387494, 25.8153961279, -77.6914895371};
test_label[1225] = '{21.1714845864};
test_output[1225] = '{51.7519025828};
############ END DEBUG ############*/
test_input[9808:9815] = '{32'h424fc6b9, 32'hc2a4d95d, 32'h41e30666, 32'h4296ef19, 32'hc26f998a, 32'h41edd00d, 32'hc217df2a, 32'h40a1aa76};
test_label[1226] = '{32'h41edd00d};
test_output[1226] = '{32'h4236f62c};
/*############ DEBUG ############
test_input[9808:9815] = '{51.9440650396, -82.4245379818, 28.3781245196, 75.4669894536, -59.899941485, 29.7265867763, -37.9679349258, 5.05205819965};
test_label[1226] = '{29.7265867763};
test_output[1226] = '{45.7404026774};
############ END DEBUG ############*/
test_input[9816:9823] = '{32'h429de2e2, 32'h42c58ab0, 32'h4116526e, 32'hc283c985, 32'hc13f461a, 32'h42bb3e26, 32'h41d66ba0, 32'h427ba461};
test_label[1227] = '{32'h429de2e2};
test_output[1227] = '{32'h419eab14};
/*############ DEBUG ############
test_input[9816:9823] = '{78.9431267698, 98.7708751601, 9.39512442035, -65.893592415, -11.9546142804, 93.6213872861, 26.8025510559, 62.9105267517};
test_label[1227] = '{78.9431267698};
test_output[1227] = '{19.8335339993};
############ END DEBUG ############*/
test_input[9824:9831] = '{32'h41d8a31f, 32'h421d83fb, 32'hc2890416, 32'h4047d5a0, 32'h423a42fe, 32'h42516829, 32'h424b3918, 32'h41e8be00};
test_label[1228] = '{32'hc2890416};
test_output[1228] = '{32'h42f21c5f};
/*############ DEBUG ############
test_input[9824:9831] = '{27.0796486938, 39.3788868474, -68.5079797854, 3.12241354847, 46.5654223177, 52.3517184232, 50.8057554442, 29.0927729485};
test_label[1228] = '{-68.5079797854};
test_output[1228] = '{121.055411534};
############ END DEBUG ############*/
test_input[9832:9839] = '{32'h419e3378, 32'hc20ef1c0, 32'h4236d14f, 32'h4299412d, 32'h42bc74fd, 32'h421a547c, 32'h4278b605, 32'h420bc7e9};
test_label[1229] = '{32'h42bc74fd};
test_output[1229] = '{32'h32c2ef1b};
/*############ DEBUG ############
test_input[9832:9839] = '{19.7751316662, -35.7360825255, 45.7044010735, 76.6272960651, 94.2284924706, 38.5825042922, 62.177753785, 34.9452239262};
test_label[1229] = '{94.2284924706};
test_output[1229] = '{2.26933050484e-08};
############ END DEBUG ############*/
test_input[9840:9847] = '{32'hc293e7e5, 32'h41c6f2b9, 32'h428f1e94, 32'hc13120cc, 32'hc126364d, 32'h41522184, 32'h42011342, 32'hc1703ee8};
test_label[1230] = '{32'h42011342};
test_output[1230] = '{32'h421d29e7};
/*############ DEBUG ############
test_input[9840:9847] = '{-73.952921256, 24.8685173574, 71.5597248919, -11.0705073611, -10.388256668, 13.1331820809, 32.2688054593, -15.0153578555};
test_label[1230] = '{32.2688054593};
test_output[1230] = '{39.2909194326};
############ END DEBUG ############*/
test_input[9848:9855] = '{32'h419ca96d, 32'hc08858f7, 32'hc288a56f, 32'hc1f433ed, 32'h4288c572, 32'hc2a533fc, 32'hbec07393, 32'hc25b27f8};
test_label[1231] = '{32'h419ca96d};
test_output[1231] = '{32'h4243362d};
/*############ DEBUG ############
test_input[9848:9855] = '{19.5827278994, -4.26085984522, -68.3231151045, -30.5253538055, 68.3856335556, -82.6015316279, -0.375881748512, -54.7890312535};
test_label[1231] = '{19.5827278994};
test_output[1231] = '{48.8029056561};
############ END DEBUG ############*/
test_input[9856:9863] = '{32'hc2b824bc, 32'h42aabc38, 32'h410a65ef, 32'hc2bf9d85, 32'hc28490ff, 32'hc05d36ae, 32'hc19dd310, 32'h42871df1};
test_label[1232] = '{32'hc19dd310};
test_output[1232] = '{32'h42d230fc};
/*############ DEBUG ############
test_input[9856:9863] = '{-92.0717501551, 85.3676181281, 8.64988629239, -95.8076553313, -66.2831984195, -3.45646247004, -19.7280577588, 67.5584816857};
test_label[1232] = '{-19.7280577588};
test_output[1232] = '{105.095675905};
############ END DEBUG ############*/
test_input[9864:9871] = '{32'hc124e1a2, 32'h4296d3af, 32'h4265f594, 32'h4219f0c5, 32'hc27ca66c, 32'h42b0bdaf, 32'hc1b45929, 32'h423dd0a5};
test_label[1233] = '{32'hc124e1a2};
test_output[1233] = '{32'h42c559e3};
/*############ DEBUG ############
test_input[9864:9871] = '{-10.3050859843, 75.4134452556, 57.4898215446, 38.4851260088, -63.1625199507, 88.3704730033, -22.5435357522, 47.4537551078};
test_label[1233] = '{-10.3050859843};
test_output[1233] = '{98.6755613472};
############ END DEBUG ############*/
test_input[9872:9879] = '{32'hc16f6004, 32'hc2ba4866, 32'hc2801e29, 32'h42834b47, 32'hc243e40f, 32'h42136cc9, 32'hc26ad1be, 32'h418d2edb};
test_label[1234] = '{32'hc26ad1be};
test_output[1234] = '{32'h42f8b426};
/*############ DEBUG ############
test_input[9872:9879] = '{-14.960941418, -93.1414011404, -64.0589029807, 65.6470263509, -48.9727122008, 36.8562368564, -58.7048255379, 17.6478786307};
test_label[1234] = '{-58.7048255379};
test_output[1234] = '{124.351851889};
############ END DEBUG ############*/
test_input[9880:9887] = '{32'hc28d8881, 32'h42acf738, 32'hc1299cb4, 32'hc2bb603d, 32'hc27d850c, 32'h425d51e9, 32'h42b0a31a, 32'h42b49871};
test_label[1235] = '{32'hc2bb603d};
test_output[1235] = '{32'h43382262};
/*############ DEBUG ############
test_input[9880:9887] = '{-70.7666055511, 86.4828460918, -10.6007579268, -93.6879672648, -63.3799286064, 55.329988539, 88.3185589785, 90.2977355638};
test_label[1235] = '{-93.6879672648};
test_output[1235] = '{184.134315162};
############ END DEBUG ############*/
test_input[9888:9895] = '{32'hc2973fa6, 32'hc2829e10, 32'h42378101, 32'h42198cdf, 32'h4232d447, 32'hc2a83121, 32'hc28920e8, 32'h410c092c};
test_label[1236] = '{32'hc2829e10};
test_output[1236] = '{32'h42dee957};
/*############ DEBUG ############
test_input[9888:9895] = '{-75.6243110825, -65.3087173561, 45.8759800576, 38.3875677955, 44.7073011713, -84.0959557159, -68.5642674217, 8.75223894504};
test_label[1236] = '{-65.3087173561};
test_output[1236] = '{111.455744468};
############ END DEBUG ############*/
test_input[9896:9903] = '{32'hc2c775b1, 32'h410f4e62, 32'hc281aee8, 32'hc22316cb, 32'h424964ad, 32'h4280a6e5, 32'h42713543, 32'h40a83973};
test_label[1237] = '{32'h424964ad};
test_output[1237] = '{32'h415fed11};
/*############ DEBUG ############
test_input[9896:9903] = '{-99.7298647825, 8.95663686268, -64.8416110342, -40.772257264, 50.3483146307, 64.3259672315, 60.3020116441, 5.25701279355};
test_label[1237] = '{50.3483146307};
test_output[1237] = '{13.9953775231};
############ END DEBUG ############*/
test_input[9904:9911] = '{32'hc20127a4, 32'hc19911e9, 32'h42147559, 32'h420e302d, 32'h42a3fe37, 32'h4237f118, 32'hc2497dfa, 32'hc287bb3b};
test_label[1238] = '{32'hc20127a4};
test_output[1238] = '{32'h42e49208};
/*############ DEBUG ############
test_input[9904:9911] = '{-32.2887099953, -19.1337443618, 37.1145965827, 35.5470471508, 81.9965097447, 45.9854445087, -50.3730230177, -67.8656838094};
test_label[1238] = '{-32.2887099953};
test_output[1238] = '{114.28521974};
############ END DEBUG ############*/
test_input[9912:9919] = '{32'hc1bd4ccb, 32'h42a96352, 32'h422affc2, 32'h4217f6c9, 32'h42bca0e7, 32'h416499ee, 32'h42046a8a, 32'h42b8a3ff};
test_label[1239] = '{32'h416499ee};
test_output[1239] = '{32'h42a04f0c};
/*############ DEBUG ############
test_input[9912:9919] = '{-23.662496087, 84.6939822054, 42.7497639622, 37.9910001181, 94.3142599544, 14.2875801976, 33.1040438575, 92.3203073597};
test_label[1239] = '{14.2875801976};
test_output[1239] = '{80.1543889729};
############ END DEBUG ############*/
test_input[9920:9927] = '{32'h424c449e, 32'hc2677983, 32'h42bb14ed, 32'hc2090a07, 32'hc22cb177, 32'hc2b5d54b, 32'h4279f250, 32'h42a2e464};
test_label[1240] = '{32'h42bb14ed};
test_output[1240] = '{32'h36bb84e9};
/*############ DEBUG ############
test_input[9920:9927] = '{51.0670081561, -57.8686639919, 93.5408695936, -34.2597923746, -43.1733038489, -90.9165879299, 62.4866315369, 81.4460740025};
test_label[1240] = '{93.5408695936};
test_output[1240] = '{5.58850706173e-06};
############ END DEBUG ############*/
test_input[9928:9935] = '{32'hc151b899, 32'hc24f9e8b, 32'hc26944da, 32'h41c3b63c, 32'h4247a54c, 32'hc11e7878, 32'hc2b0c6a6, 32'hc23eac74};
test_label[1241] = '{32'hc24f9e8b};
test_output[1241] = '{32'h42cba1eb};
/*############ DEBUG ############
test_input[9928:9935] = '{-13.1075675858, -51.9048256266, -58.3172394714, 24.4639806942, 49.9114232255, -9.9044108995, -88.3879823102, -47.6684108263};
test_label[1241] = '{-51.9048256266};
test_output[1241] = '{101.816248852};
############ END DEBUG ############*/
test_input[9936:9943] = '{32'h41f72dc8, 32'h41002020, 32'h420ac9d7, 32'hc2afe03b, 32'hc2c4f9ab, 32'h426737db, 32'hc16cd6db, 32'hc24f83e5};
test_label[1242] = '{32'hc24f83e5};
test_output[1242] = '{32'h42db5de0};
/*############ DEBUG ############
test_input[9936:9943] = '{30.8973534039, 8.00784348908, 34.6971076406, -87.9379518213, -98.4876321935, 57.8045452253, -14.8024546233, -51.8788044356};
test_label[1242] = '{-51.8788044356};
test_output[1242] = '{109.683349661};
############ END DEBUG ############*/
test_input[9944:9951] = '{32'hc216e6de, 32'hc0af04ee, 32'hc2032f46, 32'h42b85ebd, 32'h4219219c, 32'h3e87aeba, 32'hc124c939, 32'h420eb50d};
test_label[1243] = '{32'hc0af04ee};
test_output[1243] = '{32'h42c34f0c};
/*############ DEBUG ############
test_input[9944:9951] = '{-37.7254563876, -5.46935156201, -32.796164513, 92.1850340525, 38.2828200322, 0.265004931095, -10.299126525, 35.6768080752};
test_label[1243] = '{-5.46935156201};
test_output[1243] = '{97.6543856145};
############ END DEBUG ############*/
test_input[9952:9959] = '{32'h4163a6cd, 32'h42c46818, 32'hc1a1414c, 32'hc206f9c6, 32'h418842c7, 32'h425b9122, 32'h42725b1d, 32'h40802b91};
test_label[1244] = '{32'hc1a1414c};
test_output[1244] = '{32'h42ecb86b};
/*############ DEBUG ############
test_input[9952:9959] = '{14.2282230761, 98.2033056854, -20.1568825898, -33.7439201249, 17.0326052345, 54.8917322923, 60.5889790446, 4.00531829724};
test_label[1244] = '{-20.1568825898};
test_output[1244] = '{118.360188275};
############ END DEBUG ############*/
test_input[9960:9967] = '{32'h41f980c3, 32'hc282924b, 32'hc26ac4ca, 32'h42ba081b, 32'h41343cea, 32'hc2c76492, 32'hc28c3b07, 32'h4270dc98};
test_label[1245] = '{32'hc28c3b07};
test_output[1245] = '{32'h43232191};
/*############ DEBUG ############
test_input[9960:9967] = '{31.1878716189, -65.2857317987, -58.6921777089, 93.0158308364, 11.2648711783, -99.6964252916, -70.1152868938, 60.2154234875};
test_label[1245] = '{-70.1152868938};
test_output[1245] = '{163.13111773};
############ END DEBUG ############*/
test_input[9968:9975] = '{32'h429e131a, 32'h425437ae, 32'hc2688a57, 32'h411ad0e1, 32'hc237e38a, 32'hc290768f, 32'hc24e8dd9, 32'hc2425db4};
test_label[1246] = '{32'hc24e8dd9};
test_output[1246] = '{32'h4302ad03};
/*############ DEBUG ############
test_input[9968:9975] = '{79.0373050095, 53.0543737195, -58.1350993874, 9.67599575861, -45.9722047048, -72.2315562269, -51.6385222154, -48.5915051787};
test_label[1246] = '{-51.6385222154};
test_output[1246] = '{130.675827225};
############ END DEBUG ############*/
test_input[9976:9983] = '{32'h41cf4144, 32'h425002df, 32'h429a3251, 32'h426ac41a, 32'h40fd4f9b, 32'hc28c142b, 32'h4272638d, 32'h42c7696c};
test_label[1247] = '{32'h40fd4f9b};
test_output[1247] = '{32'h42b79472};
/*############ DEBUG ############
test_input[9976:9983] = '{25.906867085, 52.0028023324, 77.0982705941, 58.6915040095, 7.9159673366, -70.0393868058, 60.5972181469, 99.7059024287};
test_label[1247] = '{7.9159673366};
test_output[1247] = '{91.7899350923};
############ END DEBUG ############*/
test_input[9984:9991] = '{32'hc290f6ed, 32'hc1aea628, 32'hc1c5a099, 32'hc226d322, 32'h42aade7a, 32'h4296af85, 32'hc2ae5fd2, 32'h3f1f1a8c};
test_label[1248] = '{32'hc226d322};
test_output[1248] = '{32'h42fe4811};
/*############ DEBUG ############
test_input[9984:9991] = '{-72.482276526, -21.8311306912, -24.703417585, -41.7061842817, 85.4345282646, 75.3428112695, -87.1871495245, 0.621498818828};
test_label[1248] = '{-41.7061842817};
test_output[1248] = '{127.140753967};
############ END DEBUG ############*/
test_input[9992:9999] = '{32'h41a0f3d4, 32'h421a9c40, 32'hc06fb5e0, 32'hc23e164e, 32'h42be9323, 32'h420e2f03, 32'hc2601788, 32'hc2a08591};
test_label[1249] = '{32'h41a0f3d4};
test_output[1249] = '{32'h4296562e};
/*############ DEBUG ############
test_input[9992:9999] = '{20.1190570242, 38.6525886042, -3.74547582387, -47.5217804631, 95.2873731438, 35.545910437, -56.0229780351, -80.2608697144};
test_label[1249] = '{20.1190570242};
test_output[1249] = '{75.1683161196};
############ END DEBUG ############*/
test_input[10000:10007] = '{32'hc28a23a2, 32'hc20b6d28, 32'h429a1e90, 32'h42932f45, 32'h42b1e471, 32'h4196d973, 32'h41b57497, 32'hc1f0e986};
test_label[1250] = '{32'hc20b6d28};
test_output[1250] = '{32'h42f79b06};
/*############ DEBUG ############
test_input[10000:10007] = '{-69.0695939046, -34.8565975831, 77.0596899511, 73.5923234257, 88.9461761771, 18.8561771877, 22.6819279365, -30.114025391};
test_label[1250] = '{-34.8565975831};
test_output[1250] = '{123.802780858};
############ END DEBUG ############*/
test_input[10008:10015] = '{32'h41a6001b, 32'h424fafe9, 32'hc1ecb9c7, 32'h42b599ff, 32'hc1fe2ba7, 32'h42a1addb, 32'h4180fc97, 32'hc2960786};
test_label[1251] = '{32'hc1fe2ba7};
test_output[1251] = '{32'h42f524ef};
/*############ DEBUG ############
test_input[10008:10015] = '{20.7500512349, 51.9217853844, -29.5907113646, 90.8007716035, -31.7713146575, 80.8395633489, 16.1233347984, -75.0146957551};
test_label[1251] = '{-31.7713146575};
test_output[1251] = '{122.572133455};
############ END DEBUG ############*/
test_input[10016:10023] = '{32'h4277ec11, 32'hc260c5ce, 32'h41fe7aef, 32'h42968a2e, 32'hc26ba1e6, 32'hc1bfbf8a, 32'hc0ff8e74, 32'hc27e47b9};
test_label[1252] = '{32'h41fe7aef};
test_output[1252] = '{32'h422dd6e4};
/*############ DEBUG ############
test_input[10016:10023] = '{61.9805348357, -56.1931688258, 31.8100268139, 75.2698800975, -58.9081035087, -23.9685253999, -7.98613936698, -63.5700433976};
test_label[1252] = '{31.8100268139};
test_output[1252] = '{43.459854976};
############ END DEBUG ############*/
test_input[10024:10031] = '{32'hc2940341, 32'hc245c00a, 32'hc1f1aef6, 32'hc18b79e0, 32'h422de485, 32'h41b8e8e5, 32'hc2a9c8c4, 32'hc28c8028};
test_label[1253] = '{32'h422de485};
test_output[1253] = '{32'h30c5bfc2};
/*############ DEBUG ############
test_input[10024:10031] = '{-74.0063535148, -49.4375390053, -30.2104310604, -17.4345097144, 43.4731643843, 23.1137175367, -84.892120805, -70.2503056624};
test_label[1253] = '{43.4731643843};
test_output[1253] = '{1.43881373586e-09};
############ END DEBUG ############*/
test_input[10032:10039] = '{32'hc298d348, 32'hc276bf35, 32'hc29223a4, 32'hc2a21020, 32'h427d6f6b, 32'h42742a1a, 32'hc0ef150b, 32'hc28486d2};
test_label[1254] = '{32'hc0ef150b};
test_output[1254] = '{32'h428dd920};
/*############ DEBUG ############
test_input[10032:10039] = '{-76.4126558684, -61.6867239179, -73.0696105966, -81.0314914539, 63.3588082917, 61.0411136382, -7.4713185437, -66.2633208714};
test_label[1254] = '{-7.4713185437};
test_output[1254] = '{70.9240728139};
############ END DEBUG ############*/
test_input[10040:10047] = '{32'hc2c756d4, 32'h42acbc98, 32'hc2abd095, 32'h4225547a, 32'h424e5a2e, 32'h42c74c3f, 32'hc1d5ab95, 32'h41eaafbf};
test_label[1255] = '{32'h41eaafbf};
test_output[1255] = '{32'h428ca04f};
/*############ DEBUG ############
test_input[10040:10047] = '{-99.6695851062, 86.3683452372, -85.9073856077, 41.3324959723, 51.5880664928, 99.6489172545, -26.7087811459, 29.3358131008};
test_label[1255] = '{29.3358131008};
test_output[1255] = '{70.3131058611};
############ END DEBUG ############*/
test_input[10048:10055] = '{32'hc15246f4, 32'hc02da297, 32'hc2aa280e, 32'h42bfe6de, 32'h42be406d, 32'hc260c758, 32'hc29c0e5b, 32'hc286b763};
test_label[1256] = '{32'hc260c758};
test_output[1256] = '{32'h4318824c};
/*############ DEBUG ############
test_input[10048:10055] = '{-13.1423221707, -2.71304870982, -85.0782347299, 95.9509154557, 95.1258294601, -56.1946706005, -78.0280396756, -67.3581789473};
test_label[1256] = '{-56.1946706005};
test_output[1256] = '{152.508976516};
############ END DEBUG ############*/
test_input[10056:10063] = '{32'h42906180, 32'h42c6d729, 32'h41d195d2, 32'hc22a0b98, 32'h41a3a394, 32'h4246495a, 32'h41c83316, 32'hc2a12700};
test_label[1257] = '{32'h4246495a};
test_output[1257] = '{32'h424764f7};
/*############ DEBUG ############
test_input[10056:10063] = '{72.1904263653, 99.420233308, 26.198153607, -42.5113217845, 20.4548725323, 49.5716341066, 25.0249449258, -80.5761737242};
test_label[1257] = '{49.5716341066};
test_output[1257] = '{49.8485992014};
############ END DEBUG ############*/
test_input[10064:10071] = '{32'h42235c2b, 32'h42a9d455, 32'hc08f9732, 32'h4289d2f4, 32'h41bed55d, 32'h425bc0c2, 32'h42b6c3d3, 32'hc17b977a};
test_label[1258] = '{32'hc08f9732};
test_output[1258] = '{32'h42bfbe11};
/*############ DEBUG ############
test_input[10064:10071] = '{40.8400084532, 84.91471104, -4.48720652171, 68.9120202794, 23.8541819125, 54.9382401473, 91.382467556, -15.7244818389};
test_label[1258] = '{-4.48720652171};
test_output[1258] = '{95.871225579};
############ END DEBUG ############*/
test_input[10072:10079] = '{32'h4201e2cd, 32'h42ac31e2, 32'hc1605ff1, 32'hc27b23d1, 32'hc24139bf, 32'h4265da6d, 32'hc21c4b68, 32'h4287c6a0};
test_label[1259] = '{32'hc1605ff1};
test_output[1259] = '{32'h42c83de0};
/*############ DEBUG ############
test_input[10072:10079] = '{32.4714843911, 86.0974239228, -14.0234235927, -62.784976021, -48.3063926605, 57.4633046354, -39.0736385781, 67.8879377878};
test_label[1259] = '{-14.0234235927};
test_output[1259] = '{100.120847528};
############ END DEBUG ############*/
test_input[10080:10087] = '{32'hc2b28cf8, 32'hc2bd9cac, 32'hc2b6e972, 32'hc2a3e32c, 32'hc09fb845, 32'hc09acfce, 32'h42709031, 32'h42762b0e};
test_label[1260] = '{32'hc2bd9cac};
test_output[1260] = '{32'h431c9177};
/*############ DEBUG ############
test_input[10080:10087] = '{-89.2753294877, -94.806002757, -91.4559465386, -81.9436945533, -4.99124374706, -4.83786688951, 60.14081094, 61.542044778};
test_label[1260] = '{-94.806002757};
test_output[1260] = '{156.568220993};
############ END DEBUG ############*/
test_input[10088:10095] = '{32'h42c1049d, 32'h424c225c, 32'h40bf5c56, 32'hc179d751, 32'h422fb2a3, 32'hc274604f, 32'hc19b65ee, 32'h4262fb2e};
test_label[1261] = '{32'h4262fb2e};
test_output[1261] = '{32'h421f0e0c};
/*############ DEBUG ############
test_input[10088:10095] = '{96.5090092094, 51.0335546151, 5.98002167932, -15.6150675513, 43.9244507418, -61.0940523356, -19.4247709745, 56.745293007};
test_label[1261] = '{56.745293007};
test_output[1261] = '{39.7637162023};
############ END DEBUG ############*/
test_input[10096:10103] = '{32'h428a1847, 32'hc103edd7, 32'hc2aa632b, 32'h42b5cad0, 32'hc117876f, 32'hc18794fa, 32'h42506fd8, 32'h41ec22db};
test_label[1262] = '{32'h42506fd8};
test_output[1262] = '{32'h421b25c7};
/*############ DEBUG ############
test_input[10096:10103] = '{69.0474138842, -8.24556679126, -85.1936848012, 90.8961168089, -9.47056526101, -16.9477420522, 52.10922355, 29.5170193715};
test_label[1262] = '{52.10922355};
test_output[1262] = '{38.7868932593};
############ END DEBUG ############*/
test_input[10104:10111] = '{32'h426d4337, 32'h40916bb9, 32'hc23ffb97, 32'hc02e8dc6, 32'h4217751f, 32'hc27e6cf4, 32'h41b53b0b, 32'h42a0d31c};
test_label[1263] = '{32'h41b53b0b};
test_output[1263] = '{32'h426708b3};
/*############ DEBUG ############
test_input[10104:10111] = '{59.3156380176, 4.5443999321, -47.9956914187, -2.72740318327, 37.8643765918, -63.6064000435, 22.6538301901, 80.412324811};
test_label[1263] = '{22.6538301901};
test_output[1263] = '{57.7584946216};
############ END DEBUG ############*/
test_input[10112:10119] = '{32'hc2c6b9c7, 32'hc27b80e3, 32'h422b93ff, 32'h42803910, 32'hc1117c98, 32'hc0d97afd, 32'h4282a6f7, 32'hc296aa24};
test_label[1264] = '{32'h4282a6f7};
test_output[1264] = '{32'h3e8512f1};
/*############ DEBUG ############
test_input[10112:10119] = '{-99.3628461276, -62.8758655357, 42.8945262372, 64.1114495191, -9.09291870452, -6.79626335963, 65.3261006004, -75.3323063754};
test_label[1264] = '{65.3261006004};
test_output[1264] = '{0.259910148053};
############ END DEBUG ############*/
test_input[10120:10127] = '{32'hc0e6bebf, 32'hc2bb5691, 32'h41b96321, 32'h41c93ae4, 32'h41a075d9, 32'h42277a51, 32'hc0dd25fa, 32'hc2aced4a};
test_label[1265] = '{32'hc0e6bebf};
test_output[1265] = '{32'h42445229};
/*############ DEBUG ############
test_input[10120:10127] = '{-7.21078438227, -93.6690738756, 23.1734024643, 25.1537549171, 20.0575426049, 41.8694482277, -6.91088602376, -86.4634527747};
test_label[1265] = '{-7.21078438227};
test_output[1265] = '{49.0802326729};
############ END DEBUG ############*/
test_input[10128:10135] = '{32'h41654c9d, 32'hc2885fae, 32'h420354ba, 32'h4210fe8a, 32'h42883ca7, 32'h420ff3b8, 32'hc23e45e5, 32'hc2169fc6};
test_label[1266] = '{32'hc2885fae};
test_output[1266] = '{32'h43084e2b};
/*############ DEBUG ############
test_input[10128:10135] = '{14.3312044323, -68.1868775654, 32.8327393076, 36.2485732303, 68.1184648794, 35.9880063354, -47.5682570466, -37.6560280771};
test_label[1266] = '{-68.1868775654};
test_output[1266] = '{136.305342445};
############ END DEBUG ############*/
test_input[10136:10143] = '{32'hc156c495, 32'h42893268, 32'hc258a252, 32'h4236fa8f, 32'h42aa1622, 32'hc2022d6e, 32'h42391999, 32'hc099dd45};
test_label[1267] = '{32'h42893268};
test_output[1267] = '{32'h41838eea};
/*############ DEBUG ############
test_input[10136:10143] = '{-13.4229939884, 68.5984490469, -54.158517198, 45.744685743, 85.0432308112, -32.5443635788, 46.2749987797, -4.80826052314};
test_label[1267] = '{68.5984490469};
test_output[1267] = '{16.4447818364};
############ END DEBUG ############*/
test_input[10144:10151] = '{32'h409ee793, 32'h4222f5e6, 32'hc214e9d6, 32'h42b417e9, 32'h425f591f, 32'hc2c5c3a5, 32'h3f5b37e5, 32'h42c22dfe};
test_label[1268] = '{32'hc214e9d6};
test_output[1268] = '{32'h430651ae};
/*############ DEBUG ############
test_input[10144:10151] = '{4.96576829496, 40.740137061, -37.2283542133, 90.0466994968, 55.8370330166, -98.8821150281, 0.856321606909, 97.0898319527};
test_label[1268] = '{-37.2283542133};
test_output[1268] = '{134.319059171};
############ END DEBUG ############*/
test_input[10152:10159] = '{32'h424e908e, 32'hc2746f7e, 32'h4144f870, 32'h42c49054, 32'hbfceedda, 32'h42044231, 32'hc2bb2856, 32'hc2bf6afd};
test_label[1269] = '{32'h4144f870};
test_output[1269] = '{32'h42abf146};
/*############ DEBUG ############
test_input[10152:10159] = '{51.6411672154, -61.1088781258, 12.3106532968, 98.2818890595, -1.61663368199, 33.0646403712, -93.5787846162, -95.7089583564};
test_label[1269] = '{12.3106532968};
test_output[1269] = '{85.9712357626};
############ END DEBUG ############*/
test_input[10160:10167] = '{32'hbfb11353, 32'hc2776c76, 32'h41572e6a, 32'h412db3c9, 32'h416c2353, 32'hc0bad8fa, 32'h4213bc94, 32'h429c9fc2};
test_label[1270] = '{32'hc2776c76};
test_output[1270] = '{32'h430c2afe};
/*############ DEBUG ############
test_input[10160:10167] = '{-1.38340218573, -61.8559171203, 13.4488314989, 10.8563924466, 14.7586242334, -5.83898624101, 36.9341570394, 78.3120251496};
test_label[1270] = '{-61.8559171203};
test_output[1270] = '{140.16794227};
############ END DEBUG ############*/
test_input[10168:10175] = '{32'h423c567c, 32'hc29a31a7, 32'h41fa5014, 32'hc15fa1ca, 32'hc1a11714, 32'hc2202cfb, 32'h4292b203, 32'hc0f87ce8};
test_label[1271] = '{32'hc0f87ce8};
test_output[1271] = '{32'h42a239d1};
/*############ DEBUG ############
test_input[10168:10175] = '{47.0844559437, -77.0969767291, 31.2891004125, -13.9769994928, -20.136268187, -40.0439253683, 73.3476756542, -7.76524753683};
test_label[1271] = '{-7.76524753683};
test_output[1271] = '{81.112923191};
############ END DEBUG ############*/
test_input[10176:10183] = '{32'hc06e411d, 32'h42a22535, 32'h42a703c5, 32'h4280104e, 32'h42659f2c, 32'hc2b5d720, 32'hc2586b94, 32'h4255c6ab};
test_label[1272] = '{32'hc2b5d720};
test_output[1272] = '{32'h432e82f3};
/*############ DEBUG ############
test_input[10176:10183] = '{-3.72272416616, 81.0726735999, 83.5073624694, 64.0318471746, 57.405439727, -90.9201654898, -54.1050549025, 53.4440101512};
test_label[1272] = '{-90.9201654898};
test_output[1272] = '{174.511524387};
############ END DEBUG ############*/
test_input[10184:10191] = '{32'h4284cf2e, 32'h42a4016e, 32'h422bc738, 32'h424540a5, 32'h41701328, 32'h42bde9da, 32'h42a68b7c, 32'h42bb4b19};
test_label[1273] = '{32'h41701328};
test_output[1273] = '{32'h42a061c2};
/*############ DEBUG ############
test_input[10184:10191] = '{66.4046499484, 82.0027958956, 42.9445500683, 49.3131285617, 15.0046771074, 94.9567414213, 83.2724307626, 93.6466747729};
test_label[1273] = '{15.0046771074};
test_output[1273] = '{80.1909338537};
############ END DEBUG ############*/
test_input[10192:10199] = '{32'h42c0880e, 32'hc1a79c7d, 32'h42680a65, 32'hc25fc3dd, 32'h3e8d5993, 32'h42bf8415, 32'h41805c4a, 32'hc293676d};
test_label[1274] = '{32'h3e8d5993};
test_output[1274] = '{32'h42c0ebef};
/*############ DEBUG ############
test_input[10192:10199] = '{96.2657290355, -20.9514102704, 58.0101492463, -55.9412709982, 0.276074016993, 95.7579708169, 16.0450621734, -73.7020012214};
test_label[1274] = '{0.276074016993};
test_output[1274] = '{96.4608100276};
############ END DEBUG ############*/
test_input[10200:10207] = '{32'h42c3b652, 32'h42b95aad, 32'hc23eb477, 32'h424b3f9f, 32'hc2332182, 32'hc2799249, 32'hc1ac5969, 32'h408f4336};
test_label[1275] = '{32'hc2332182};
test_output[1275] = '{32'h430ea4fa};
/*############ DEBUG ############
test_input[10200:10207] = '{97.8560978553, 92.6771000658, -47.6762336161, 50.8121294775, -44.7827218989, -62.3928561972, -21.5436568687, 4.47695468664};
test_label[1275] = '{-44.7827218989};
test_output[1275] = '{142.644437594};
############ END DEBUG ############*/
test_input[10208:10215] = '{32'h41aef55d, 32'h42058c9c, 32'hc191bffe, 32'h4296e9c3, 32'hc284e6be, 32'hc1b6e2be, 32'hc12c21e3, 32'h42b81250};
test_label[1276] = '{32'hc284e6be};
test_output[1276] = '{32'h431e7c87};
/*############ DEBUG ############
test_input[10208:10215] = '{21.8698054041, 33.3873157156, -18.2187459662, 75.4565648098, -66.450667742, -22.8607138715, -10.7582729669, 92.0357681159};
test_label[1276] = '{-66.450667742};
test_output[1276] = '{158.486435921};
############ END DEBUG ############*/
test_input[10216:10223] = '{32'hc2063943, 32'hc2b1abc0, 32'hc226fae5, 32'hc27d1134, 32'hc26578bb, 32'hc2272da5, 32'h42a985f8, 32'hc23451eb};
test_label[1277] = '{32'hc2063943};
test_output[1277] = '{32'h42eca29a};
/*############ DEBUG ############
test_input[10216:10223] = '{-33.5559178354, -88.8354511967, -41.7450148472, -63.266801165, -57.3679010567, -41.7945751686, 84.7616607503, -45.0799990832};
test_label[1277] = '{-33.5559178354};
test_output[1277] = '{118.317578586};
############ END DEBUG ############*/
test_input[10224:10231] = '{32'h426fcc72, 32'h427abaeb, 32'hc2c69f9a, 32'h42458f20, 32'h4280d045, 32'hc2c7c4a1, 32'h42b97743, 32'hc07e9b74};
test_label[1278] = '{32'h4280d045};
test_output[1278] = '{32'h41e29bf6};
/*############ DEBUG ############
test_input[10224:10231] = '{59.9496530503, 62.6825389412, -99.3117203351, 49.3897702423, 64.4067762929, -99.8840430951, 92.7329297575, -3.97823809606};
test_label[1278] = '{64.4067762929};
test_output[1278] = '{28.3261534646};
############ END DEBUG ############*/
test_input[10232:10239] = '{32'h41c4b9de, 32'hc21535c3, 32'hc192cb89, 32'hc266a5fa, 32'h4240b400, 32'h421b183c, 32'h42889eb3, 32'hc2884032};
test_label[1279] = '{32'hc266a5fa};
test_output[1279] = '{32'h42fbf1b0};
/*############ DEBUG ############
test_input[10232:10239] = '{24.590755912, -37.3025023979, -18.3493818994, -57.6620847832, 48.175781244, 38.7736650998, 68.3099627421, -68.1253821399};
test_label[1279] = '{-57.6620847832};
test_output[1279] = '{125.972047527};
############ END DEBUG ############*/
test_input[10240:10247] = '{32'h41e4f9a8, 32'h42c6331d, 32'h428e1b64, 32'h4263107c, 32'h42a6085f, 32'h42aaedfb, 32'h42b276bc, 32'hc1c03020};
test_label[1280] = '{32'h42aaedfb};
test_output[1280] = '{32'h415a2948};
/*############ DEBUG ############
test_input[10240:10247] = '{28.6219021747, 99.0998294934, 71.0534936317, 56.7660984114, 83.0163526744, 85.4648044126, 89.2319013282, -24.0234989936};
test_label[1280] = '{85.4648044126};
test_output[1280] = '{13.6350781907};
############ END DEBUG ############*/
test_input[10248:10255] = '{32'hc29b4a0a, 32'hc2c6b6a8, 32'h418a85b8, 32'h427e42eb, 32'h42c0783d, 32'h42b39f2a, 32'h4252120c, 32'h42a5620e};
test_label[1281] = '{32'h427e42eb};
test_output[1281] = '{32'h4202af38};
/*############ DEBUG ############
test_input[10248:10255] = '{-77.6446046773, -99.3567495065, 17.3152920991, 63.5653479272, 96.2348369843, 89.8108663632, 52.5176231666, 82.6915141409};
test_label[1281] = '{63.5653479272};
test_output[1281] = '{32.6711112557};
############ END DEBUG ############*/
test_input[10256:10263] = '{32'hc29abd56, 32'hc26c3548, 32'h42784eae, 32'hc1cd2956, 32'h4150e741, 32'hc266f9ef, 32'hc2077db3, 32'hc28f623a};
test_label[1282] = '{32'h4150e741};
test_output[1282] = '{32'h424414de};
/*############ DEBUG ############
test_input[10256:10263] = '{-77.3697975321, -59.052031812, 62.0768352697, -25.6451828243, 13.0564580474, -57.7440744861, -33.8727542805, -71.691846378};
test_label[1282] = '{13.0564580474};
test_output[1282] = '{49.0203772223};
############ END DEBUG ############*/
test_input[10264:10271] = '{32'hc18539e4, 32'hc2ac4fdc, 32'h422cd277, 32'hc23e280f, 32'hc20accfc, 32'h42874339, 32'h4290a7e3, 32'hc2b03cc6};
test_label[1283] = '{32'hc20accfc};
test_output[1283] = '{32'h42d61307};
/*############ DEBUG ############
test_input[10264:10271] = '{-16.6532669632, -86.1559740562, 43.205533805, -47.5391194409, -34.7001792863, 67.6312914407, 72.3279024365, -88.1186955457};
test_label[1283] = '{-34.7001792863};
test_output[1283] = '{107.037166484};
############ END DEBUG ############*/
test_input[10272:10279] = '{32'h41e23bbf, 32'h42a11946, 32'hc20333df, 32'hc2bdc775, 32'h422bfc62, 32'hc23c1164, 32'h41fc0a22, 32'hc0903775};
test_label[1284] = '{32'h41fc0a22};
test_output[1284] = '{32'h42442d7b};
/*############ DEBUG ############
test_input[10272:10279] = '{28.279172991, 80.5493629356, -32.8006557795, -94.8895616204, 42.9964667241, -47.016981442, 31.5049485831, -4.50676955064};
test_label[1284] = '{31.5049485831};
test_output[1284] = '{49.0444143525};
############ END DEBUG ############*/
test_input[10280:10287] = '{32'h42946734, 32'h428afd55, 32'h421f4dda, 32'h4293cab9, 32'hc172990a, 32'h42b23be6, 32'hc1839fa2, 32'h423fcd2b};
test_label[1285] = '{32'hc172990a};
test_output[1285] = '{32'h42d08f07};
/*############ DEBUG ############
test_input[10280:10287] = '{74.2015714173, 69.4947855895, 39.8260278841, 73.8959402642, -15.162362652, 89.1169893692, -16.4529449903, 47.9503575357};
test_label[1285] = '{-15.162362652};
test_output[1285] = '{104.279352602};
############ END DEBUG ############*/
test_input[10288:10295] = '{32'h42757531, 32'h412403dd, 32'h41a833b8, 32'hc25712df, 32'h42b443e6, 32'hc2abd317, 32'h4281dc8d, 32'h42bbeca2};
test_label[1286] = '{32'h4281dc8d};
test_output[1286] = '{32'h41e86c56};
/*############ DEBUG ############
test_input[10288:10295] = '{61.3644443736, 10.2509430168, 21.0252524192, -53.7684306641, 90.1326170391, -85.9122881554, 64.9307628631, 93.9621743123};
test_label[1286] = '{64.9307628631};
test_output[1286] = '{29.0528981765};
############ END DEBUG ############*/
test_input[10296:10303] = '{32'h41df0c87, 32'h4234878d, 32'h42a33a8a, 32'hc21d1a49, 32'hc2adb6e5, 32'hc2892e25, 32'hc2bbea51, 32'hc1ce77f6};
test_label[1287] = '{32'hc1ce77f6};
test_output[1287] = '{32'h42d6d888};
/*############ DEBUG ############
test_input[10296:10303] = '{27.8811163909, 45.132375208, 81.6143345895, -39.2756701431, -86.8572159036, -68.5901245769, -93.9576521844, -25.8085753028};
test_label[1287] = '{-25.8085753028};
test_output[1287] = '{107.422909892};
############ END DEBUG ############*/
test_input[10304:10311] = '{32'h4284d58e, 32'h41c951cb, 32'h427d7786, 32'hc29daecd, 32'h42bc9923, 32'h42a35586, 32'hc1fec03d, 32'hc2b0d147};
test_label[1288] = '{32'hc1fec03d};
test_output[1288] = '{32'h42fc4933};
/*############ DEBUG ############
test_input[10304:10311] = '{66.4171023975, 25.164937374, 63.3667211819, -78.8414049476, 94.2990966992, 81.6670407825, -31.8438654041, -88.4087447332};
test_label[1288] = '{-31.8438654041};
test_output[1288] = '{126.142965369};
############ END DEBUG ############*/
test_input[10312:10319] = '{32'h42067fee, 32'hc243500b, 32'h42a6899c, 32'h429675c2, 32'h42a496d3, 32'h426b3e0d, 32'h42c623cd, 32'h42877446};
test_label[1289] = '{32'h42067fee};
test_output[1289] = '{32'h4282e3d6};
/*############ DEBUG ############
test_input[10312:10319] = '{33.6249313489, -48.8281675474, 83.2687664693, 75.2299989587, 82.2945750169, 58.8105948911, 99.069923268, 67.7270962396};
test_label[1289] = '{33.6249313489};
test_output[1289] = '{65.4449921083};
############ END DEBUG ############*/
test_input[10320:10327] = '{32'hc21b542d, 32'hc1fa3bf0, 32'hc1b25d7b, 32'h421ac59a, 32'h42882598, 32'hc1e35a2d, 32'h41b511f6, 32'h41eff4be};
test_label[1290] = '{32'hc21b542d};
test_output[1290] = '{32'h42d5cfae};
/*############ DEBUG ############
test_input[10320:10327] = '{-38.8322013347, -31.279266147, -22.2956454803, 38.6929708314, 68.0734241616, -28.419031567, 22.6337692383, 29.9945037847};
test_label[1290] = '{-38.8322013347};
test_output[1290] = '{106.905625496};
############ END DEBUG ############*/
test_input[10328:10335] = '{32'h3f06695f, 32'h42a43496, 32'hc2b4f34c, 32'h42bab9d4, 32'hc2b5fb52, 32'h426d9754, 32'h42ba83c0, 32'hc2bca646};
test_label[1291] = '{32'hc2b4f34c};
test_output[1291] = '{32'h43387ad9};
/*############ DEBUG ############
test_input[10328:10335] = '{0.525045362238, 82.1027040113, -90.4751863415, 93.3629429708, -90.9908618571, 59.3977813344, 93.257322185, -94.3247532323};
test_label[1291] = '{-90.4751863415};
test_output[1291] = '{184.479866698};
############ END DEBUG ############*/
test_input[10336:10343] = '{32'h411712e8, 32'h423b8c4c, 32'h4205a590, 32'hc17ca486, 32'h42374566, 32'h42b9cbf4, 32'h41608c7e, 32'hc2ab565f};
test_label[1292] = '{32'hc17ca486};
test_output[1292] = '{32'h42d96085};
/*############ DEBUG ############
test_input[10336:10343] = '{9.44211598727, 46.8870075938, 33.4116835215, -15.7901669315, 45.8177709739, 92.8983441834, 14.0343001863, -85.6686902854};
test_label[1292] = '{-15.7901669315};
test_output[1292] = '{108.688511115};
############ END DEBUG ############*/
test_input[10344:10351] = '{32'h42a4d1c8, 32'hc29b66b2, 32'h42b0b371, 32'h428977f7, 32'h424e143e, 32'hc274e4f6, 32'hc22a92fa, 32'hc1e523c8};
test_label[1293] = '{32'h42a4d1c8};
test_output[1293] = '{32'h40be300c};
/*############ DEBUG ############
test_input[10344:10351] = '{82.4097295179, -77.7005735713, 88.3504679547, 68.734305563, 51.5197682433, -61.2235934891, -42.6435300452, -28.6424709009};
test_label[1293] = '{82.4097295179};
test_output[1293] = '{5.94336507399};
############ END DEBUG ############*/
test_input[10352:10359] = '{32'hc15ba504, 32'hc26a3dda, 32'h413ee129, 32'hc1ef57f8, 32'h41baffe0, 32'h42a7d279, 32'h427145e5, 32'h40eb753e};
test_label[1294] = '{32'h42a7d279};
test_output[1294] = '{32'h2e7979e0};
/*############ DEBUG ############
test_input[10352:10359] = '{-13.7277873544, -58.5604038074, 11.9299708692, -29.9179530477, 23.3749390883, 83.911075938, 60.3182570111, 7.35806162765};
test_label[1294] = '{83.911075938};
test_output[1294] = '{5.67242919319e-11};
############ END DEBUG ############*/
test_input[10360:10367] = '{32'h42ac85a5, 32'h42337cc8, 32'hc26fc99f, 32'hc26c47fa, 32'h413061b6, 32'h4293d8fc, 32'h42830fca, 32'h424cf52c};
test_label[1295] = '{32'h42ac85a5};
test_output[1295] = '{32'h36932eb4};
/*############ DEBUG ############
test_input[10360:10367] = '{86.2610250561, 44.8718571576, -59.9468943479, -59.0702902326, 11.0238556324, 73.9237941541, 65.5308363972, 51.2394268118};
test_label[1295] = '{86.2610250561};
test_output[1295] = '{4.38637828132e-06};
############ END DEBUG ############*/
test_input[10368:10375] = '{32'h426e8739, 32'hc26df948, 32'hc29a9a33, 32'hc2083d89, 32'hc2b87319, 32'hc28c59ba, 32'hc278d863, 32'h428a0282};
test_label[1296] = '{32'hc29a9a33};
test_output[1296] = '{32'h43124e60};
/*############ DEBUG ############
test_input[10368:10375] = '{59.6320526208, -59.4934388356, -77.3011732364, -34.060094284, -92.2248007551, -70.1752472706, -62.2113166856, 69.0048973316};
test_label[1296] = '{-77.3011732364};
test_output[1296] = '{146.306155566};
############ END DEBUG ############*/
test_input[10376:10383] = '{32'hc1340527, 32'hc0a85d65, 32'hc2a45b60, 32'hc238363b, 32'h41413ff8, 32'hc2a93ce7, 32'hc2828687, 32'hc1afb5df};
test_label[1297] = '{32'hc1340527};
test_output[1297] = '{32'h41baa28f};
/*############ DEBUG ############
test_input[10376:10383] = '{-11.2512577676, -5.26140083357, -82.1784694083, -46.0529586997, 12.0781173435, -84.6189493333, -65.2627456907, -21.963803848};
test_label[1297] = '{-11.2512577676};
test_output[1297] = '{23.3293751406};
############ END DEBUG ############*/
test_input[10384:10391] = '{32'h425776ad, 32'h4230648c, 32'h42c41ef7, 32'hc21a4774, 32'hc2943aa0, 32'hc2abcaf9, 32'h42ad4a88, 32'h41a730f8};
test_label[1298] = '{32'hc21a4774};
test_output[1298] = '{32'h4308a159};
/*############ DEBUG ############
test_input[10384:10391] = '{53.8658940773, 44.0981908001, 98.0604769842, -38.5697768878, -74.1145002645, -85.8964293031, 86.6455715525, 20.8989097168};
test_label[1298] = '{-38.5697768878};
test_output[1298] = '{136.630264902};
############ END DEBUG ############*/
test_input[10392:10399] = '{32'h42c25667, 32'h4212756f, 32'h42548b77, 32'h4216b997, 32'h4077df84, 32'hc2ab26e1, 32'h41609f50, 32'h428bda80};
test_label[1299] = '{32'h4212756f};
test_output[1299] = '{32'h4272375f};
/*############ DEBUG ############
test_input[10392:10399] = '{97.1687517514, 36.6146797112, 53.1361959536, 37.6812413423, 3.873017402, -85.5759350799, 14.0388949837, 69.9267585447};
test_label[1299] = '{36.6146797112};
test_output[1299] = '{60.5540720402};
############ END DEBUG ############*/
test_input[10400:10407] = '{32'hc21cb0fb, 32'h42600094, 32'h4217562c, 32'hc2c6b8cd, 32'h41011511, 32'hc2877f60, 32'hc29094e7, 32'hc2ad0f41};
test_label[1300] = '{32'hc29094e7};
test_output[1300] = '{32'h43004a99};
/*############ DEBUG ############
test_input[10400:10407] = '{-39.1728330546, 56.0005662572, 37.8341522406, -99.3609424889, 8.06764358178, -67.7487779379, -72.2908269102, -86.5297927339};
test_label[1300] = '{-72.2908269102};
test_output[1300] = '{128.29139318};
############ END DEBUG ############*/
test_input[10408:10415] = '{32'hc289f5d1, 32'hc25ff2d6, 32'h419731b1, 32'h425fafa9, 32'h41fec2f3, 32'hc0335597, 32'hc24670f1, 32'h423687c9};
test_label[1301] = '{32'h423687c9};
test_output[1301] = '{32'h41249fa4};
/*############ DEBUG ############
test_input[10408:10415] = '{-68.9801076391, -55.9871429461, 18.8992626214, 55.9215435261, 31.8451907357, -2.80209906328, -49.6102953858, 45.6326026337};
test_label[1301] = '{45.6326026337};
test_output[1301] = '{10.288974899};
############ END DEBUG ############*/
test_input[10416:10423] = '{32'hc285c17c, 32'h427a3378, 32'h428565ef, 32'h42a5c3de, 32'h429667c5, 32'hc237922b, 32'h420f2002, 32'h42b30072};
test_label[1302] = '{32'h428565ef};
test_output[1302] = '{32'h41b66cc7};
/*############ DEBUG ############
test_input[10416:10423] = '{-66.8778958546, 62.5502617519, 66.6990886729, 82.8825502919, 75.202678187, -45.8927428908, 35.7812559093, 89.500867455};
test_label[1302] = '{66.6990886729};
test_output[1302] = '{22.803114184};
############ END DEBUG ############*/
test_input[10424:10431] = '{32'hc18167d5, 32'h415feb59, 32'hc1e5c654, 32'hc12d7480, 32'hc2997c54, 32'h4251fd44, 32'h421ccfa6, 32'hc216e76a};
test_label[1303] = '{32'h421ccfa6};
test_output[1303] = '{32'h4154b678};
/*############ DEBUG ############
test_input[10424:10431] = '{-16.1756991463, 13.9949579069, -28.7218402162, -10.8409420118, -76.7428291915, 52.4973303103, 39.202783496, -37.7259918345};
test_label[1303] = '{39.202783496};
test_output[1303] = '{13.2945484979};
############ END DEBUG ############*/
test_input[10432:10439] = '{32'hc2bb432a, 32'h42157c5c, 32'h4054cd24, 32'h416b86da, 32'hc2a3917f, 32'h40a8f452, 32'hc2b2969e, 32'h42289894};
test_label[1304] = '{32'h4054cd24};
test_output[1304] = '{32'h421b5457};
/*############ DEBUG ############
test_input[10432:10439] = '{-93.6311800864, 37.3714448651, 3.32502070763, 14.7204226706, -81.7841690872, 5.2798241021, -89.2941729746, 42.1490034987};
test_label[1304] = '{3.32502070763};
test_output[1304] = '{38.8323640914};
############ END DEBUG ############*/
test_input[10440:10447] = '{32'hc297a4ff, 32'hc2b555f1, 32'h42612c8f, 32'h41afe8b0, 32'h41444807, 32'hc283bb3e, 32'hc2964b6e, 32'h427461a9};
test_label[1305] = '{32'hc2964b6e};
test_output[1305] = '{32'h4308403a};
/*############ DEBUG ############
test_input[10440:10447] = '{-75.8222588589, -90.6678547318, 56.2935136103, 21.9886161028, 12.267584584, -65.8657104653, -75.1473251002, 61.0953730906};
test_label[1305] = '{-75.1473251002};
test_output[1305] = '{136.250879094};
############ END DEBUG ############*/
test_input[10448:10455] = '{32'hc2af6693, 32'h41b7c994, 32'hc1a1af74, 32'h4238be73, 32'hc2b84f7d, 32'hc24eebfc, 32'hc2a5f9c6, 32'hc2ab5b70};
test_label[1306] = '{32'hc1a1af74};
test_output[1306] = '{32'h4284cb17};
/*############ DEBUG ############
test_input[10448:10455] = '{-87.7003409574, 22.9734259603, -20.2106702115, 46.185986882, -92.1552519061, -51.7304552726, -82.9878421641, -85.6785854237};
test_label[1306] = '{-20.2106702115};
test_output[1306] = '{66.3966570935};
############ END DEBUG ############*/
test_input[10456:10463] = '{32'h3ff894f6, 32'h42af8cc6, 32'h42a92939, 32'hc186e9ed, 32'h41e84127, 32'h42c26cdb, 32'h42c491cf, 32'h420a21ed};
test_label[1307] = '{32'h3ff894f6};
test_output[1307] = '{32'h42c14634};
/*############ DEBUG ############
test_input[10456:10463] = '{1.94204590863, 87.7749458571, 84.5805158445, -16.8642218854, 29.0318127104, 97.2126065783, 98.2847844416, 34.5331294777};
test_label[1307] = '{1.94204590863};
test_output[1307] = '{96.637116157};
############ END DEBUG ############*/
test_input[10464:10471] = '{32'h41ab9c01, 32'hc2b01365, 32'h4265d553, 32'h42a79f43, 32'h42040765, 32'hc28d2829, 32'h41febf70, 32'h41497228};
test_label[1308] = '{32'hc2b01365};
test_output[1308] = '{32'h432bd954};
/*############ DEBUG ############
test_input[10464:10471] = '{21.4511733261, -88.0378763752, 57.4583227409, 83.8110585638, 33.0072208765, -70.5784373535, 31.8434746119, 12.5903705634};
test_label[1308] = '{-88.0378763752};
test_output[1308] = '{171.848934939};
############ END DEBUG ############*/
test_input[10472:10479] = '{32'hc277117e, 32'h42c6b8a8, 32'hc24e4c32, 32'h42b9b4c3, 32'h4251dfcd, 32'h415668d8, 32'hc29f9e0e, 32'hc287f375};
test_label[1309] = '{32'h4251dfcd};
test_output[1309] = '{32'h423b930a};
/*############ DEBUG ############
test_input[10472:10479] = '{-61.7670818084, 99.3606593566, -51.5744088593, 92.8530528551, 52.4685573105, 13.4005963789, -79.8087006548, -67.975501606};
test_label[1309] = '{52.4685573105};
test_output[1309] = '{46.8935929809};
############ END DEBUG ############*/
test_input[10480:10487] = '{32'hc2813853, 32'h42af9d64, 32'hc2b306ad, 32'h427cea56, 32'h4297a227, 32'h425c7e5c, 32'h429f58e2, 32'hc23fc565};
test_label[1310] = '{32'h427cea56};
test_output[1310] = '{32'h41c4a182};
/*############ DEBUG ############
test_input[10480:10487] = '{-64.6100105153, 87.8074036409, -89.5130410509, 63.228842262, 75.8167046457, 55.1233964634, 79.6736013619, -47.9427666409};
test_label[1310] = '{63.228842262};
test_output[1310] = '{24.578860986};
############ END DEBUG ############*/
test_input[10488:10495] = '{32'h428a52bb, 32'hc1abe543, 32'h41cc3b74, 32'h4245216f, 32'hc2284870, 32'h42a4ea5e, 32'hc251122d, 32'hc20598d3};
test_label[1311] = '{32'hc2284870};
test_output[1311] = '{32'h42f90e96};
/*############ DEBUG ############
test_input[10488:10495] = '{69.1615811991, -21.4869449588, 25.5290306904, 49.2826518189, -42.0707379894, 82.4577502483, -52.2677493451, -33.3992405207};
test_label[1311] = '{-42.0707379894};
test_output[1311] = '{124.528489919};
############ END DEBUG ############*/
test_input[10496:10503] = '{32'h42bc7a62, 32'hc21a109e, 32'h423f6d65, 32'h41be3c97, 32'hc22a4330, 32'hc25a133d, 32'hc2a55182, 32'h42a2f99e};
test_label[1312] = '{32'hc25a133d};
test_output[1312] = '{32'h4314c201};
/*############ DEBUG ############
test_input[10496:10503] = '{94.2390321848, -38.5162285411, 47.8568321357, 23.7795857562, -42.5656138042, -54.5187858735, -82.6591916387, 81.4875322176};
test_label[1312] = '{-54.5187858735};
test_output[1312] = '{148.757820956};
############ END DEBUG ############*/
test_input[10504:10511] = '{32'hc22782e2, 32'h425840d5, 32'hc2a224be, 32'hc2bd9752, 32'hc2a21f94, 32'h41b0eecc, 32'hc2b56477, 32'hc285d475};
test_label[1313] = '{32'hc2bd9752};
test_output[1313] = '{32'h4314dbdf};
/*############ DEBUG ############
test_input[10504:10511] = '{-41.8778161398, 54.0633140804, -81.0717595247, -94.7955510878, -81.0616785492, 22.1166009794, -90.6962189422, -66.9149537681};
test_label[1313] = '{-94.7955510878};
test_output[1313] = '{148.858865168};
############ END DEBUG ############*/
test_input[10512:10519] = '{32'hc1c7fefa, 32'h4295731f, 32'hc28196c0, 32'hc13c9160, 32'h42584bf8, 32'h4229f6b6, 32'h42a7ecc2, 32'h41eb4ef5};
test_label[1314] = '{32'h41eb4ef5};
test_output[1314] = '{32'h425a3224};
/*############ DEBUG ############
test_input[10512:10519] = '{-24.9994999011, 74.7248426464, -64.7944362855, -11.7854918942, 54.0741900521, 42.4909293334, 83.9624205084, 29.413553638};
test_label[1314] = '{29.413553638};
test_output[1314] = '{54.5489641787};
############ END DEBUG ############*/
test_input[10520:10527] = '{32'h410314cb, 32'h41d56571, 32'h423634ec, 32'hc296492f, 32'hc2063756, 32'h417a7821, 32'hc2b85330, 32'hc108055f};
test_label[1315] = '{32'hc296492f};
test_output[1315] = '{32'h42f163a5};
/*############ DEBUG ############
test_input[10520:10527] = '{8.19257618067, 26.674532132, 45.5516821997, -75.142935441, -33.5540377969, 15.6543281051, -92.1624737365, -8.5013112846};
test_label[1315] = '{-75.142935441};
test_output[1315] = '{120.694617647};
############ END DEBUG ############*/
test_input[10528:10535] = '{32'hc2950503, 32'h40a97996, 32'h42c1a6d8, 32'h42a61b97, 32'h4266cb94, 32'hc2275209, 32'hc285a44d, 32'hc2a943b4};
test_label[1316] = '{32'h42a61b97};
test_output[1316] = '{32'h415c5a0a};
/*############ DEBUG ############
test_input[10528:10535] = '{-74.5097911387, 5.29609222978, 96.8258667955, 83.0538852721, 57.6988086436, -41.830113522, -66.8209033982, -84.6322349643};
test_label[1316] = '{83.0538852721};
test_output[1316] = '{13.771982568};
############ END DEBUG ############*/
test_input[10536:10543] = '{32'h42374f61, 32'hc103f5d2, 32'hc1ee6437, 32'h41deedb2, 32'h4180977e, 32'h418ee76f, 32'hc0940de8, 32'hc223f311};
test_label[1317] = '{32'hc223f311};
test_output[1317] = '{32'h42ada139};
/*############ DEBUG ############
test_input[10536:10543] = '{45.8275172888, -8.24751439624, -29.7989323163, 27.8660630553, 16.0739698779, 17.8630045071, -4.62669743425, -40.9873713934};
test_label[1317] = '{-40.9873713934};
test_output[1317] = '{86.814888698};
############ END DEBUG ############*/
test_input[10544:10551] = '{32'hc23565b6, 32'h41b9eb1e, 32'hc2959370, 32'h42516210, 32'h41b3a4b6, 32'h42a37554, 32'h429b04e2, 32'hc2b9e25c};
test_label[1318] = '{32'hc2959370};
test_output[1318] = '{32'h431c881f};
/*############ DEBUG ############
test_input[10544:10551] = '{-45.3493270464, 23.2398025812, -74.7879641812, 52.3457642845, 22.4554246044, 81.729156166, 77.5095385949, -92.9421086271};
test_label[1318] = '{-74.7879641812};
test_output[1318] = '{156.531717554};
############ END DEBUG ############*/
test_input[10552:10559] = '{32'h4292b6da, 32'h3ed7e5bf, 32'hc199e209, 32'h42059871, 32'hc18247eb, 32'hc178af26, 32'h4250a0c6, 32'h4292079b};
test_label[1319] = '{32'h4250a0c6};
test_output[1319] = '{32'h41ade4c7};
/*############ DEBUG ############
test_input[10552:10559] = '{73.3571290698, 0.421674700758, -19.2353678372, 33.3988698858, -16.2851166199, -15.5427607235, 52.1570066352, 73.0148580703};
test_label[1319] = '{52.1570066352};
test_output[1319] = '{21.7367068696};
############ END DEBUG ############*/
test_input[10560:10567] = '{32'hc2726dfe, 32'hc128b37a, 32'h4209a26e, 32'hc19dd737, 32'h4293f45f, 32'h427b8bad, 32'h428ac39f, 32'hc2c6d3fe};
test_label[1320] = '{32'hc19dd737};
test_output[1320] = '{32'h42bb6f54};
/*############ DEBUG ############
test_input[10560:10567] = '{-60.607412848, -10.5438171905, 34.4086233258, -19.7300858218, 73.9772883056, 62.8864016383, 69.3820754754, -99.4140501782};
test_label[1320] = '{-19.7300858218};
test_output[1320] = '{93.7174386315};
############ END DEBUG ############*/
test_input[10568:10575] = '{32'hc1626baf, 32'hc1d80735, 32'hc289b284, 32'h4252f61e, 32'hc217fab8, 32'hc2637593, 32'hc249615e, 32'hc2c3d05b};
test_label[1321] = '{32'hc1d80735};
test_output[1321] = '{32'h429f7cdc};
/*############ DEBUG ############
test_input[10568:10575] = '{-14.1512900442, -27.0035196179, -68.8486615879, 52.7403489031, -37.9948434208, -56.8648176058, -50.34508425, -97.9069408333};
test_label[1321] = '{-27.0035196179};
test_output[1321] = '{79.743868521};
############ END DEBUG ############*/
test_input[10576:10583] = '{32'hc22a1cf7, 32'hc2986e16, 32'h42c7139d, 32'h42adb5d1, 32'h422b13a2, 32'hc293ee66, 32'h42a9650f, 32'h42722de9};
test_label[1322] = '{32'h42adb5d1};
test_output[1322] = '{32'h414aee67};
/*############ DEBUG ############
test_input[10576:10583] = '{-42.5282859343, -76.2150136859, 99.5383074296, 86.8551071846, 42.7691720993, -73.9656198292, 84.6973828789, 60.5448357855};
test_label[1322] = '{86.8551071846};
test_output[1322] = '{12.6832037064};
############ END DEBUG ############*/
test_input[10584:10591] = '{32'hc2802b8a, 32'h416471fc, 32'hc25000a1, 32'hc2b6cf54, 32'h41f97a63, 32'hc2a0eef6, 32'hc2beec45, 32'h421758af};
test_label[1323] = '{32'hc25000a1};
test_output[1323] = '{32'h42b3ad51};
/*############ DEBUG ############
test_input[10584:10591] = '{-64.0850397076, 14.2778281577, -52.0006130088, -91.4049404816, 31.1847591643, -80.4667241312, -95.4614629086, 37.8366039454};
test_label[1323] = '{-52.0006130088};
test_output[1323] = '{89.8385077579};
############ END DEBUG ############*/
test_input[10592:10599] = '{32'h428094ca, 32'hc2293c0e, 32'h4144bb2f, 32'h41e68745, 32'h42aac123, 32'h4292650d, 32'h429b115f, 32'h4207a33d};
test_label[1324] = '{32'hc2293c0e};
test_output[1324] = '{32'h42ff5f5e};
/*############ DEBUG ############
test_input[10592:10599] = '{64.2906010973, -42.3086472644, 12.2956993542, 28.8160493832, 85.3772224543, 73.1973674291, 77.5339254578, 33.9094113998};
test_label[1324] = '{-42.3086472644};
test_output[1324] = '{127.686267146};
############ END DEBUG ############*/
test_input[10600:10607] = '{32'h42ab4de6, 32'h42b95187, 32'hc2a3f8c0, 32'h4210301b, 32'hc2c38d70, 32'h42425e50, 32'hc286c48c, 32'hc2410493};
test_label[1325] = '{32'hc2c38d70};
test_output[1325] = '{32'h433e6fb7};
/*############ DEBUG ############
test_input[10600:10607] = '{85.6521483668, 92.6592322294, -81.9858370743, 36.0469798048, -97.7762432, 48.5921012492, -67.3838798458, -48.2544653071};
test_label[1325] = '{-97.7762432};
test_output[1325] = '{190.436380465};
############ END DEBUG ############*/
test_input[10608:10615] = '{32'h427aa278, 32'h428fd049, 32'h42c42ec1, 32'h41f2f15a, 32'hc159bed9, 32'h422d515a, 32'hc00c7d6b, 32'hc2627c94};
test_label[1326] = '{32'hc2627c94};
test_output[1326] = '{32'h431ab686};
/*############ DEBUG ############
test_input[10608:10615] = '{62.6586595688, 71.9068034041, 98.0913172938, 30.3678483008, -13.6090932456, 43.3294431383, -2.19515479433, -56.6216579171};
test_label[1326] = '{-56.6216579171};
test_output[1326] = '{154.712975211};
############ END DEBUG ############*/
test_input[10616:10623] = '{32'h4298943d, 32'h4295e926, 32'hc2210035, 32'h4289ea7a, 32'hc2b401f2, 32'h3fc22a8c, 32'h42978ed3, 32'hc195ba4b};
test_label[1327] = '{32'h42978ed3};
test_output[1327] = '{32'h3f911339};
/*############ DEBUG ############
test_input[10616:10623] = '{76.2895279252, 74.9553690315, -40.2502026875, 68.9579623003, -90.0037991291, 1.51692340754, 75.7789523784, -18.7159636854};
test_label[1327] = '{75.7789523784};
test_output[1327] = '{1.13339909157};
############ END DEBUG ############*/
test_input[10624:10631] = '{32'h427b33e3, 32'hc19cf63b, 32'h4031a9ec, 32'h42755345, 32'hc241ad3c, 32'hc28a2539, 32'h421f3175, 32'h402b2453};
test_label[1328] = '{32'h42755345};
test_output[1328] = '{32'h3fd6953a};
/*############ DEBUG ############
test_input[10624:10631] = '{62.8006724899, -19.6202295283, 2.77599617145, 61.3313176984, -48.4191734807, -69.0726972932, 39.798297592, 2.67409197462};
test_label[1328] = '{61.3313176984};
test_output[1328] = '{1.67642902658};
############ END DEBUG ############*/
test_input[10632:10639] = '{32'hc231f092, 32'hc0df536c, 32'h41d11a93, 32'hc196009b, 32'hc298f16e, 32'h4228022f, 32'h4235d4dc, 32'h41e5ccb9};
test_label[1329] = '{32'hc196009b};
test_output[1329] = '{32'h42807a7e};
/*############ DEBUG ############
test_input[10632:10639] = '{-44.4849315937, -6.97893353642, 26.1379761112, -18.750295852, -76.4715406486, 42.00213257, 45.4578695161, 28.7249617693};
test_label[1329] = '{-18.750295852};
test_output[1329] = '{64.2392415553};
############ END DEBUG ############*/
test_input[10640:10647] = '{32'hc264191d, 32'hc17bdfcb, 32'h41f5b783, 32'hc2aba2c3, 32'h41a03fb1, 32'h429187f2, 32'hc0f8a728, 32'hc2926fc4};
test_label[1330] = '{32'hc2aba2c3};
test_output[1330] = '{32'h431e955a};
/*############ DEBUG ############
test_input[10640:10647] = '{-57.0245252378, -15.7421368455, 30.7146046901, -85.8178948955, 20.0310992228, 72.7655166665, -7.77040477076, -73.2182960395};
test_label[1330] = '{-85.8178948955};
test_output[1330] = '{158.583411562};
############ END DEBUG ############*/
test_input[10648:10655] = '{32'h42933e27, 32'h4208cddd, 32'hc1afdd38, 32'h425bfba3, 32'hc2a5ad13, 32'h3ea32f81, 32'hc2811751, 32'h428296e5};
test_label[1331] = '{32'h4208cddd};
test_output[1331] = '{32'h421daeb1};
/*############ DEBUG ############
test_input[10648:10655] = '{73.6213946258, 34.2010392653, -21.9830173198, 54.9957380009, -82.8380326249, 0.318721800272, -64.5455402151, 65.2947153355};
test_label[1331] = '{34.2010392653};
test_output[1331] = '{39.4205973136};
############ END DEBUG ############*/
test_input[10656:10663] = '{32'hc1b86156, 32'hc23d97a4, 32'h41758ff1, 32'hc1f0880f, 32'hc2bcd7ea, 32'hc256dedd, 32'hc12ce38f, 32'h420190e5};
test_label[1332] = '{32'hc256dedd};
test_output[1332] = '{32'h42ac37e1};
/*############ DEBUG ############
test_input[10656:10663] = '{-23.0475270218, -47.398086211, 15.3476423527, -30.0664349795, -94.4217087968, -53.7176402205, -10.8055564042, 32.3915001784};
test_label[1332] = '{-53.7176402205};
test_output[1332] = '{86.1091404385};
############ END DEBUG ############*/
test_input[10664:10671] = '{32'h4268e6c9, 32'hc2ba5254, 32'hc2517031, 32'hc2055440, 32'hc2b4bfee, 32'hc2b23e8e, 32'hc15ca4f1, 32'h42bd4e5d};
test_label[1333] = '{32'hc2055440};
test_output[1333] = '{32'h42fff87d};
/*############ DEBUG ############
test_input[10664:10671] = '{58.2253753233, -93.1607996873, -52.359563417, -33.3322739991, -90.3748646617, -89.1221735788, -13.7902684838, 94.6530557711};
test_label[1333] = '{-33.3322739991};
test_output[1333] = '{127.98532977};
############ END DEBUG ############*/
test_input[10672:10679] = '{32'hc2a1fa85, 32'h429e4df1, 32'hc1ff3d7f, 32'hc241111c, 32'hc282f9a5, 32'hc26af7b7, 32'hc16806db, 32'h41eda91e};
test_label[1334] = '{32'hc282f9a5};
test_output[1334] = '{32'h4310a3cb};
/*############ DEBUG ############
test_input[10672:10679] = '{-80.9892930125, 79.1522313798, -31.9050267053, -48.2667069616, -65.4875878682, -58.7419081975, -14.5016734148, 29.7075760968};
test_label[1334] = '{-65.4875878682};
test_output[1334] = '{144.639819248};
############ END DEBUG ############*/
test_input[10680:10687] = '{32'hc2c6459a, 32'h42a55bb8, 32'h42a33f5f, 32'h424b3131, 32'hc1d5cf6d, 32'h416a2fd6, 32'h42a032c3, 32'h42a37568};
test_label[1335] = '{32'hc1d5cf6d};
test_output[1335] = '{32'h42dbff8b};
/*############ DEBUG ############
test_input[10680:10687] = '{-99.1359403207, 82.6791396576, 81.6237726644, 50.7980388412, -26.7262822884, 14.636679016, 80.0991417762, 81.7293064015};
test_label[1335] = '{-26.7262822884};
test_output[1335] = '{109.999104721};
############ END DEBUG ############*/
test_input[10688:10695] = '{32'h40e2222a, 32'hc2c5698b, 32'h428ec13c, 32'hc2a1d474, 32'hc220a4ab, 32'hc00322f6, 32'h41b792f4, 32'hc28436b1};
test_label[1336] = '{32'h40e2222a};
test_output[1336] = '{32'h42809f1a};
/*############ DEBUG ############
test_input[10688:10695] = '{7.06667056814, -98.7061392509, 71.3774146886, -80.9149502514, -40.1608074765, -2.04900883373, 22.9467549263, -66.1068173658};
test_label[1336] = '{7.06667056814};
test_output[1336] = '{64.3107441204};
############ END DEBUG ############*/
test_input[10696:10703] = '{32'hc0c3c099, 32'h42bce47d, 32'hc1034d48, 32'h42bd1645, 32'hc10c4335, 32'h41423075, 32'hc178eea6, 32'h42c26a56};
test_label[1337] = '{32'hc10c4335};
test_output[1337] = '{32'h42d4329b};
/*############ DEBUG ############
test_input[10696:10703] = '{-6.11726024506, 94.4462646902, -8.20636704012, 94.5434941531, -8.76640791304, 12.1368301804, -15.5582638231, 97.2076871922};
test_label[1337] = '{-8.76640791304};
test_output[1337] = '{106.098838166};
############ END DEBUG ############*/
test_input[10704:10711] = '{32'h4296f8be, 32'hc1eafb31, 32'h3f0dff47, 32'hc2619808, 32'h42c0205a, 32'hc207baef, 32'h42b8d5dd, 32'h422850a7};
test_label[1338] = '{32'h42b8d5dd};
test_output[1338] = '{32'h406af5eb};
/*############ DEBUG ############
test_input[10704:10711] = '{75.4858267083, -29.372651259, 0.554676463929, -56.3984682895, 96.0631889178, -33.9325539493, 92.4177030729, 42.0787635374};
test_label[1338] = '{92.4177030729};
test_output[1338] = '{3.67125955401};
############ END DEBUG ############*/
test_input[10712:10719] = '{32'h4287b0c7, 32'h42c00325, 32'h425775f8, 32'h42634106, 32'hc20814aa, 32'hc27db80a, 32'h413373dd, 32'hc2298cbf};
test_label[1339] = '{32'h4287b0c7};
test_output[1339] = '{32'h41e14977};
/*############ DEBUG ############
test_input[10712:10719] = '{67.845267599, 96.0061383064, 53.8652024525, 56.8134986164, -34.0201779994, -63.4297239778, 11.2157872956, -42.3874473377};
test_label[1339] = '{67.845267599};
test_output[1339] = '{28.1608707074};
############ END DEBUG ############*/
test_input[10720:10727] = '{32'hc2733879, 32'h3ffa6d25, 32'h42857d03, 32'hc23c0283, 32'hc2a9f8a6, 32'h41ee700a, 32'h4267bb6d, 32'hc2aedc41};
test_label[1340] = '{32'h41ee700a};
test_output[1340] = '{32'h4213c227};
/*############ DEBUG ############
test_input[10720:10727] = '{-60.8051502221, 1.95645586774, 66.7441609501, -47.0024516332, -84.9856419089, 29.8047062421, 57.933032829, -87.4301798213};
test_label[1340] = '{29.8047062421};
test_output[1340] = '{36.9396037619};
############ END DEBUG ############*/
test_input[10728:10735] = '{32'h42359cf7, 32'h4253efe1, 32'hc0b794f2, 32'hc260ba55, 32'hc2c379cf, 32'hc1bd02cb, 32'hc222a325, 32'hc1ed16c6};
test_label[1341] = '{32'h42359cf7};
test_output[1341] = '{32'h40f29b7e};
/*############ DEBUG ############
test_input[10728:10735] = '{45.4032853374, 52.9842564933, -5.73693165767, -56.1819650095, -97.7379092287, -23.6263645213, -40.6593205374, -29.6361189564};
test_label[1341] = '{45.4032853374};
test_output[1341] = '{7.58148109151};
############ END DEBUG ############*/
test_input[10736:10743] = '{32'h42b2893e, 32'hc101695c, 32'h4232437f, 32'hc2478fab, 32'h42af7e91, 32'hc28c2ac8, 32'hc227b45b, 32'h41d613b2};
test_label[1342] = '{32'h4232437f};
test_output[1342] = '{32'h42339960};
/*############ DEBUG ############
test_input[10736:10743] = '{89.2680534833, -8.08822237472, 44.5659135147, -49.8903010855, 87.7472011213, -70.0835551918, -41.9261269626, 26.7596171993};
test_label[1342] = '{44.5659135147};
test_output[1342] = '{44.8997815265};
############ END DEBUG ############*/
test_input[10744:10751] = '{32'h42104da4, 32'hc29c50cf, 32'h429185cc, 32'h41ef371f, 32'hc1e13b0d, 32'hc20fcf3f, 32'hc2854a55, 32'hc20d2e17};
test_label[1343] = '{32'hc20d2e17};
test_output[1343] = '{32'h42d81cd7};
/*############ DEBUG ############
test_input[10744:10751] = '{36.075820003, -78.1578260285, 72.7613194305, 29.9019152256, -28.1538337818, -35.9523889054, -66.6451782105, -35.2950103959};
test_label[1343] = '{-35.2950103959};
test_output[1343] = '{108.056329826};
############ END DEBUG ############*/
test_input[10752:10759] = '{32'h428f06b4, 32'h42401c2d, 32'hc26a8f1b, 32'hc1a49c9e, 32'h428e5c6e, 32'hc2816784, 32'h418ef83a, 32'h42c06eb7};
test_label[1344] = '{32'h42c06eb7};
test_output[1344] = '{32'h2e0d2080};
/*############ DEBUG ############
test_input[10752:10759] = '{71.5130923093, 48.0275151663, -58.6397516828, -20.5764735059, 71.1805266773, -64.702178007, 17.8712041123, 96.2162420852};
test_label[1344] = '{96.2162420852};
test_output[1344] = '{3.20885540367e-11};
############ END DEBUG ############*/
test_input[10760:10767] = '{32'hc22df62d, 32'hc29627fc, 32'h41894307, 32'h4234cc1c, 32'h428b7c59, 32'h42b97743, 32'h41220c49, 32'h419e28d9};
test_label[1345] = '{32'hc22df62d};
test_output[1345] = '{32'h4308392d};
/*############ DEBUG ############
test_input[10760:10767] = '{-43.490407815, -75.0780917347, 17.1577290424, 45.1993271292, 69.7428667488, 92.7329351838, 10.1279988534, 19.7699448446};
test_label[1345] = '{-43.490407815};
test_output[1345] = '{136.223342999};
############ END DEBUG ############*/
test_input[10768:10775] = '{32'h4299fd6b, 32'h42388667, 32'h421100ab, 32'hc18599e8, 32'hc2154c7b, 32'h4155eccb, 32'hc24aae8c, 32'h427f2aac};
test_label[1346] = '{32'h421100ab};
test_output[1346] = '{32'h4222fa2c};
/*############ DEBUG ############
test_input[10768:10775] = '{76.9949598712, 46.1312540554, 36.2506513791, -16.7001494747, -37.3246864343, 13.3703105976, -50.6704544748, 63.7916707823};
test_label[1346] = '{36.2506513791};
test_output[1346] = '{40.7443103367};
############ END DEBUG ############*/
test_input[10776:10783] = '{32'h428029e4, 32'h41252c15, 32'hc0c5fd00, 32'h4251fe49, 32'hc12f33e7, 32'hc2a03fdd, 32'h41070609, 32'hc2a0936d};
test_label[1347] = '{32'hc2a0936d};
test_output[1347] = '{32'h43105ea9};
/*############ DEBUG ############
test_input[10776:10783] = '{64.0818172637, 10.3232617631, -6.18713360241, 52.4983270148, -10.9501715313, -80.1247313069, 8.43897387508, -80.2879441138};
test_label[1347] = '{-80.2879441138};
test_output[1347] = '{144.369770696};
############ END DEBUG ############*/
test_input[10784:10791] = '{32'hc222836e, 32'h42bcd64e, 32'h41ea8208, 32'h423cff41, 32'h40ca275d, 32'h424a08ef, 32'h4253063b, 32'hc14d24a1};
test_label[1348] = '{32'h41ea8208};
test_output[1348] = '{32'h428235cc};
/*############ DEBUG ############
test_input[10784:10791] = '{-40.628347901, 94.4185626029, 29.3134912262, 47.2492700853, 6.31730504122, 50.5087237279, 52.7560827113, -12.8214422014};
test_label[1348] = '{29.3134912262};
test_output[1348] = '{65.1050713767};
############ END DEBUG ############*/
test_input[10792:10799] = '{32'h42902f08, 32'hc23d98e2, 32'hc2151ba8, 32'hc2b68c88, 32'h42726ccc, 32'hc22dc153, 32'hc2b84ac8, 32'hc2c7c357};
test_label[1349] = '{32'hc2b84ac8};
test_output[1349] = '{32'h43243ce9};
/*############ DEBUG ############
test_input[10792:10799] = '{72.0918559189, -47.3993015123, -37.2770075426, -91.2744735793, 60.6062465403, -43.4387935767, -92.1460567141, -99.8815194026};
test_label[1349] = '{-92.1460567141};
test_output[1349] = '{164.23792291};
############ END DEBUG ############*/
test_input[10800:10807] = '{32'hc2c2765a, 32'h42c05825, 32'h42ba19fe, 32'h42b2daf7, 32'hc1d2da9c, 32'hc0b0d527, 32'hc27dde6e, 32'h425762dd};
test_label[1350] = '{32'h42c05825};
test_output[1350] = '{32'h3d355d0e};
/*############ DEBUG ############
test_input[10800:10807] = '{-97.231154555, 96.1721592526, 93.0507676754, 89.4276640534, -26.3567432005, -5.52601935275, -63.467217451, 53.8465479071};
test_label[1350] = '{96.1721592526};
test_output[1350] = '{0.0442781966303};
############ END DEBUG ############*/
test_input[10808:10815] = '{32'h4178ee04, 32'hc2a12f82, 32'h41c1ad5c, 32'h42b06d05, 32'hc2acf136, 32'h42c25d29, 32'hc04e6794, 32'h42b223b0};
test_label[1351] = '{32'hc2a12f82};
test_output[1351] = '{32'h4331c671};
/*############ DEBUG ############
test_input[10808:10815] = '{15.5581091169, -80.5927877592, 24.2096483343, 88.2129294762, -86.471115746, 97.1819535078, -3.22507190162, 89.0697054118};
test_label[1351] = '{-80.5927877592};
test_output[1351] = '{177.775168312};
############ END DEBUG ############*/
test_input[10816:10823] = '{32'h41f76b4b, 32'h42c42dd9, 32'hc1897f3a, 32'hc1d31b45, 32'h42b9733c, 32'hc2c1e864, 32'hbf825740, 32'hc1a5ca35};
test_label[1352] = '{32'hc1897f3a};
test_output[1352] = '{32'h42e6900b};
/*############ DEBUG ############
test_input[10816:10823] = '{30.9273896819, 98.0895425691, -17.1871222891, -26.3883159599, 92.725068459, -96.9538846896, -1.01828764907, -20.7237335423};
test_label[1352] = '{-17.1871222891};
test_output[1352] = '{115.281333862};
############ END DEBUG ############*/
test_input[10824:10831] = '{32'h418147e0, 32'h4215f587, 32'hc2507505, 32'hc1c85311, 32'hc170bd03, 32'h424f36c3, 32'hc1b2e763, 32'hc0b147d2};
test_label[1353] = '{32'hc1b2e763};
test_output[1353] = '{32'h4294553a};
/*############ DEBUG ############
test_input[10824:10831] = '{16.1600947858, 37.4897719013, -52.1142779159, -25.0405606165, -15.0461451516, 51.8034770974, -22.3629820844, -5.54001699842};
test_label[1353] = '{-22.3629820844};
test_output[1353] = '{74.1664597895};
############ END DEBUG ############*/
test_input[10832:10839] = '{32'h4148a5f3, 32'h428f73bf, 32'hc1a40a5e, 32'h4256d8da, 32'h42a5d294, 32'hc2a92951, 32'h4233b899, 32'h41d32cad};
test_label[1354] = '{32'h41d32cad};
test_output[1354] = '{32'h42620ed5};
/*############ DEBUG ############
test_input[10832:10839] = '{12.5405146148, 71.7260666564, -20.5050623025, 53.7117678138, 82.9112870219, -84.580693412, 44.9302715783, 26.3968146367};
test_label[1354] = '{26.3968146367};
test_output[1354] = '{56.5144862629};
############ END DEBUG ############*/
test_input[10840:10847] = '{32'hc21d5571, 32'hc0a411c9, 32'hc2822df0, 32'hc15afc82, 32'hc2846c55, 32'hc293bc07, 32'hc26c75ba, 32'h42415745};
test_label[1355] = '{32'hc2822df0};
test_output[1355] = '{32'h42e2d992};
/*############ DEBUG ############
test_input[10840:10847] = '{-39.3334404278, -5.12717119481, -65.0897182922, -13.6866478152, -66.2115894712, -73.8672388935, -59.1149667063, 48.3352233885};
test_label[1355] = '{-65.0897182922};
test_output[1355] = '{113.424941681};
############ END DEBUG ############*/
test_input[10848:10855] = '{32'hc299de3a, 32'h410b4d6e, 32'h4244c191, 32'hc2794e2d, 32'h425f6285, 32'hc2872b12, 32'h42b4a5c9, 32'h42c4778e};
test_label[1356] = '{32'hc2794e2d};
test_output[1356] = '{32'h43208f6b};
/*############ DEBUG ############
test_input[10848:10855] = '{-76.934039873, 8.70640375908, 49.189029852, -62.3263452644, 55.8462094408, -67.5841197162, 90.3237955345, 98.2335085545};
test_label[1356] = '{-62.3263452644};
test_output[1356] = '{160.560220911};
############ END DEBUG ############*/
test_input[10856:10863] = '{32'hc1cb13f2, 32'h42926158, 32'h425452d7, 32'h41bacac2, 32'hc2722963, 32'hc181881e, 32'hc2a4e5e5, 32'h420e1d09};
test_label[1357] = '{32'hc2722963};
test_output[1357] = '{32'h4305bb04};
/*############ DEBUG ############
test_input[10856:10863] = '{-25.3847387755, 73.190121885, 53.0808968528, 23.3490028524, -60.5404153859, -16.1914626561, -82.4490126017, 35.5283534632};
test_label[1357] = '{-60.5404153859};
test_output[1357] = '{133.730537273};
############ END DEBUG ############*/
test_input[10864:10871] = '{32'hc213416a, 32'hc240d148, 32'h40b1ae0b, 32'hc11f1214, 32'hc146c40e, 32'h425b9988, 32'hc22c8427, 32'hc29f9332};
test_label[1358] = '{32'hc240d148};
test_output[1358] = '{32'h42ce3568};
/*############ DEBUG ############
test_input[10864:10871] = '{-36.8138818356, -48.2043775604, 5.55249531538, -9.94191386543, -12.422864928, 54.8999314215, -43.1290567869, -79.7874938831};
test_label[1358] = '{-48.2043775604};
test_output[1358] = '{103.104308982};
############ END DEBUG ############*/
test_input[10872:10879] = '{32'hc2983e04, 32'hc1cbb665, 32'h42765e55, 32'h40d79380, 32'h41c727e6, 32'h41e40c9e, 32'h41d1acc3, 32'h428e8e9f};
test_label[1359] = '{32'h40d79380};
test_output[1359] = '{32'h4281156f};
/*############ DEBUG ############
test_input[10872:10879] = '{-76.1211270852, -25.4640603935, 61.5921193607, 6.73675525949, 24.8944816275, 28.5061614954, 26.2093559336, 71.2785557369};
test_label[1359] = '{6.73675525949};
test_output[1359] = '{64.5418625958};
############ END DEBUG ############*/
test_input[10880:10887] = '{32'h426bab1d, 32'h410e9f4a, 32'h41d152ed, 32'hc19f8801, 32'hc1fcfd8c, 32'hc24d0f0e, 32'hc13a5874, 32'h3f2dcfcc};
test_label[1360] = '{32'hc24d0f0e};
test_output[1360] = '{32'h42dc5d16};
/*############ DEBUG ############
test_input[10880:10887] = '{58.9171029245, 8.91388855583, 26.1654911205, -19.9414073325, -31.6238019612, -51.2647033867, -11.6465949957, 0.678951964992};
test_label[1360] = '{-51.2647033867};
test_output[1360] = '{110.181806311};
############ END DEBUG ############*/
test_input[10888:10895] = '{32'h4288b946, 32'hc2725afa, 32'h41b80f86, 32'hc28e217e, 32'h423fd5c9, 32'h426a8169, 32'h42406096, 32'hc2aa7dbd};
test_label[1361] = '{32'h426a8169};
test_output[1361] = '{32'h411bc4c7};
/*############ DEBUG ############
test_input[10888:10895] = '{68.3618593696, -60.5888431842, 23.007579153, -71.0654144758, 47.9587734852, 58.6263770181, 48.0943211936, -85.2455839402};
test_label[1361] = '{58.6263770181};
test_output[1361] = '{9.73554149986};
############ END DEBUG ############*/
test_input[10896:10903] = '{32'h42767671, 32'hc2383bc1, 32'h42bc9356, 32'h424ead5d, 32'h417d21c2, 32'h41f78966, 32'h420d52a4, 32'hc2a2c49a};
test_label[1362] = '{32'h42bc9356};
test_output[1362] = '{32'h27ec0000};
/*############ DEBUG ############
test_input[10896:10903] = '{61.6156635871, -46.0583540629, 94.2877638351, 51.6692991551, 15.8207413171, 30.9420899957, 35.3307052974, -81.3839866924};
test_label[1362] = '{94.2877638351};
test_output[1362] = '{6.55031584529e-15};
############ END DEBUG ############*/
test_input[10904:10911] = '{32'h42425061, 32'hc22115ad, 32'hc208e416, 32'h3fc02ec9, 32'h4111a117, 32'hc2b7bb92, 32'h42aa4509, 32'hc2785ad4};
test_label[1363] = '{32'hc22115ad};
test_output[1363] = '{32'h42facfe0};
/*############ DEBUG ############
test_input[10904:10911] = '{48.5784957958, -40.2711677978, -34.2227420399, 1.50142782084, 9.10182866892, -91.8663486991, 85.1348349532, -62.0886985408};
test_label[1363] = '{-40.2711677978};
test_output[1363] = '{125.406002751};
############ END DEBUG ############*/
test_input[10912:10919] = '{32'hc2a7b039, 32'h42858a9f, 32'hc2094e80, 32'h4294dd5b, 32'h424693cc, 32'hc262c69f, 32'hc2772c0a, 32'hc1cfc78a};
test_label[1364] = '{32'hc2a7b039};
test_output[1364] = '{32'h431e46e8};
/*############ DEBUG ############
test_input[10912:10919] = '{-83.8441811181, 66.7707466594, -34.3266604032, 74.4323313807, 49.6443325789, -56.6939667568, -61.7930056066, -25.9724314985};
test_label[1364] = '{-83.8441811181};
test_output[1364] = '{158.276982949};
############ END DEBUG ############*/
test_input[10920:10927] = '{32'hc2996c82, 32'h423aee3f, 32'h425210d8, 32'hc204865f, 32'h42a9a62e, 32'hc2154360, 32'h4279453b, 32'h4211623d};
test_label[1365] = '{32'h4279453b};
test_output[1365] = '{32'h41b40e44};
/*############ DEBUG ############
test_input[10920:10927] = '{-76.7119269604, 46.7326612701, 52.5164499214, -33.1312217387, 84.8245721376, -37.3157974155, 62.3176059738, 36.3459356522};
test_label[1365] = '{62.3176059738};
test_output[1365] = '{22.506966164};
############ END DEBUG ############*/
test_input[10928:10935] = '{32'hc2c0b477, 32'h42a90e59, 32'hc2995c81, 32'h414cddcb, 32'hc229c773, 32'hc1ef89e1, 32'hc27affcb, 32'hc2379d3b};
test_label[1366] = '{32'hc2c0b477};
test_output[1366] = '{32'h4334e168};
/*############ DEBUG ############
test_input[10928:10935] = '{-96.3524667404, 84.5280249867, -76.6806729958, 12.8041489203, -42.4447728553, -29.9423239474, -62.7497967567, -45.9035450612};
test_label[1366] = '{-96.3524667404};
test_output[1366] = '{180.880491727};
############ END DEBUG ############*/
test_input[10936:10943] = '{32'hc263bbf2, 32'h42871929, 32'hc1af591c, 32'hc2818686, 32'h41ed23c4, 32'h425628c0, 32'h428c8d88, 32'hc23a8530};
test_label[1367] = '{32'hc263bbf2};
test_output[1367] = '{32'h42fe8bf0};
/*############ DEBUG ############
test_input[10936:10943] = '{-56.933540223, 67.5491410952, -21.9185101196, -64.762737657, 29.6424638607, 53.5397944955, 70.2764315716, -46.6300658795};
test_label[1367] = '{-56.933540223};
test_output[1367] = '{127.273318634};
############ END DEBUG ############*/
test_input[10944:10951] = '{32'h418b5bdd, 32'h41c5e95b, 32'h429cdc7d, 32'h42a0b034, 32'h42968ed1, 32'h3f59e100, 32'h428677c0, 32'hc2a0fcd0};
test_label[1368] = '{32'hc2a0fcd0};
test_output[1368] = '{32'h4320fb26};
/*############ DEBUG ############
test_input[10944:10951] = '{17.4198558093, 24.7389437938, 78.4306397675, 80.3441485797, 75.2789357513, 0.851089448384, 67.2338843157, -80.4937736408};
test_label[1368] = '{-80.4937736408};
test_output[1368] = '{160.981049193};
############ END DEBUG ############*/
test_input[10952:10959] = '{32'hc25da1fb, 32'hc1f6546f, 32'hc276071e, 32'hc0c22a19, 32'hc2207b5c, 32'h41d55be3, 32'hc0689f56, 32'hc17c7a8f};
test_label[1369] = '{32'hc1f6546f};
test_output[1369] = '{32'h4265d829};
/*############ DEBUG ############
test_input[10952:10959] = '{-55.408182308, -30.7912272921, -61.5069508456, -6.06763898421, -40.1204676949, 26.669866253, -3.63472498431, -15.7799219021};
test_label[1369] = '{-30.7912272921};
test_output[1369] = '{57.4610935452};
############ END DEBUG ############*/
test_input[10960:10967] = '{32'h419e3d59, 32'hc20b269b, 32'hc22817f1, 32'h4225c85b, 32'hc2c3d295, 32'hc04891df, 32'hc0eb0be1, 32'h420ee502};
test_label[1370] = '{32'hc2c3d295};
test_output[1370] = '{32'h430b5c38};
/*############ DEBUG ############
test_input[10960:10967] = '{19.7799549146, -34.7877014858, -42.0233787967, 41.4456590006, -97.911295873, -3.13390332527, -7.34520017837, 35.7236388404};
test_label[1370] = '{-97.911295873};
test_output[1370] = '{139.360222621};
############ END DEBUG ############*/
test_input[10968:10975] = '{32'hc21161fc, 32'hc28363b1, 32'h4163301d, 32'h41431f7e, 32'h42a4f344, 32'hc1c6639b, 32'h42b24d50, 32'h421babcf};
test_label[1371] = '{32'h4163301d};
test_output[1371] = '{32'h4295e7f2};
/*############ DEBUG ############
test_input[10968:10975] = '{-36.3456867682, -65.6947075642, 14.1992460099, 12.1951888157, 82.4751268059, -24.7986363972, 89.1510004471, 38.9177832841};
test_label[1371] = '{14.1992460099};
test_output[1371] = '{74.9530146133};
############ END DEBUG ############*/
test_input[10976:10983] = '{32'hc09c9fbb, 32'hc2b4edee, 32'h416a125c, 32'h42005472, 32'hc2be614b, 32'h424a5734, 32'hc1ee91b5, 32'hc1da3d1b};
test_label[1372] = '{32'h416a125c};
test_output[1372] = '{32'h420fd29d};
/*############ DEBUG ############
test_input[10976:10983] = '{-4.89449849416, -90.4647066421, 14.6294824069, 32.0824646549, -95.1900229233, 50.5851597198, -29.8211453641, -27.2798371869};
test_label[1372] = '{14.6294824069};
test_output[1372] = '{35.9556773221};
############ END DEBUG ############*/
test_input[10984:10991] = '{32'h4282ddf9, 32'h420104eb, 32'h41567d5a, 32'hc2870645, 32'h42085acc, 32'hc260a8ac, 32'hc26181f1, 32'h424dae2f};
test_label[1373] = '{32'h424dae2f};
test_output[1373] = '{32'h41603709};
/*############ DEBUG ############
test_input[10984:10991] = '{65.4335366528, 32.2548019412, 13.4056036671, -67.5122417263, 34.0886706109, -56.1647186457, -56.3768973849, 51.4201012923};
test_label[1373] = '{51.4201012923};
test_output[1373] = '{14.013436181};
############ END DEBUG ############*/
test_input[10992:10999] = '{32'h414257cd, 32'hc257c1dd, 32'h42c0143e, 32'h42aaa39a, 32'h42b32738, 32'h40931f87, 32'hc27b505d, 32'h42985369};
test_label[1374] = '{32'h42aaa39a};
test_output[1374] = '{32'h412b8b9b};
/*############ DEBUG ############
test_input[10992:10999] = '{12.146435704, -53.9393205236, 96.0395362503, 85.3195340475, 89.576601625, 4.5975987796, -62.8284807279, 76.1629071119};
test_label[1374] = '{85.3195340475};
test_output[1374] = '{10.7215832634};
############ END DEBUG ############*/
test_input[11000:11007] = '{32'h4221616a, 32'hbfdcaa40, 32'h42bb3fc8, 32'h42a20b01, 32'hc283f8b8, 32'h4278c702, 32'hc2a23203, 32'h3f79ee14};
test_label[1375] = '{32'hbfdcaa40};
test_output[1375] = '{32'h42beb271};
/*############ DEBUG ############
test_input[11000:11007] = '{40.3451320439, -1.72394564549, 93.624569281, 81.0214918803, -65.98577534, 62.1943451064, -81.0976773668, 0.976289011604};
test_label[1375] = '{-1.72394564549};
test_output[1375] = '{95.3485182882};
############ END DEBUG ############*/
test_input[11008:11015] = '{32'h411a066d, 32'h42a66adc, 32'h42b15bfc, 32'h416d4b5b, 32'h428ed041, 32'h429b6711, 32'hc27b83dd, 32'hc2bcc38c};
test_label[1376] = '{32'h42a66adc};
test_output[1376] = '{32'h40af3490};
/*############ DEBUG ############
test_input[11008:11015] = '{9.62656918585, 83.2087065001, 88.6796573007, 14.8308969825, 71.4067482522, 77.7012992985, -62.8787739847, -94.3819273162};
test_label[1376] = '{83.2087065001};
test_output[1376] = '{5.47516623178};
############ END DEBUG ############*/
test_input[11016:11023] = '{32'h422b22e6, 32'hc29ecd62, 32'hc220567d, 32'h42a815ac, 32'hc19b4763, 32'hc127551b, 32'hc2871572, 32'h4282d2ce};
test_label[1377] = '{32'h4282d2ce};
test_output[1377] = '{32'h41950b76};
/*############ DEBUG ############
test_input[11016:11023] = '{42.7840793307, -79.4011378222, -40.0844607805, 84.0423259173, -19.4098577204, -10.4582773298, -67.5418820375, 65.411728941};
test_label[1377] = '{65.411728941};
test_output[1377] = '{18.6305969844};
############ END DEBUG ############*/
test_input[11024:11031] = '{32'h41ed050d, 32'hc28450f0, 32'hc2243b73, 32'hc254340f, 32'h427c717d, 32'hc2bc49c5, 32'hc0fc94e2, 32'hc2b4ab0d};
test_label[1378] = '{32'hc0fc94e2};
test_output[1378] = '{32'h428e020d};
/*############ DEBUG ############
test_input[11024:11031] = '{29.6274670008, -66.1580797013, -41.05805745, -53.0508396492, 63.1108289349, -94.1440827224, -7.8931741492, -90.334086802};
test_label[1378] = '{-7.8931741492};
test_output[1378] = '{71.0040030841};
############ END DEBUG ############*/
test_input[11032:11039] = '{32'h40b99d19, 32'hc230223b, 32'hc289cef2, 32'hc1a5a38e, 32'h41d9be4a, 32'hc21f7841, 32'hc2aeca20, 32'hc2a43cdb};
test_label[1379] = '{32'hc289cef2};
test_output[1379] = '{32'h42c03e85};
/*############ DEBUG ############
test_input[11032:11039] = '{5.80042696848, -44.0334267852, -68.9041926467, -20.7048604651, 27.217914942, -39.8674341538, -87.3947756557, -82.1188568371};
test_label[1379] = '{-68.9041926467};
test_output[1379] = '{96.1221075892};
############ END DEBUG ############*/
test_input[11040:11047] = '{32'hc2809882, 32'hc25e8d2b, 32'hc2b0c5c6, 32'hc1ec8e7d, 32'h4256a532, 32'h427e50a9, 32'h41b21fb4, 32'hc22e4b04};
test_label[1380] = '{32'hc2809882};
test_output[1380] = '{32'h42ffc0dd};
/*############ DEBUG ############
test_input[11040:11047] = '{-64.2978671352, -55.6378607941, -88.3862796388, -29.5695734557, 53.6613218846, 63.578771575, 22.2654799899, -43.5732563046};
test_label[1380] = '{-64.2978671352};
test_output[1380] = '{127.876688016};
############ END DEBUG ############*/
test_input[11048:11055] = '{32'h4271c10e, 32'hc162e922, 32'h41bd45e9, 32'h428d26c2, 32'h4205ba1b, 32'h4160a6f6, 32'h4279bc12, 32'h40bbfc0f};
test_label[1381] = '{32'hc162e922};
test_output[1381] = '{32'h42a98412};
/*############ DEBUG ############
test_input[11048:11055] = '{60.4385291034, -14.1819173741, 23.6591352139, 70.5757006589, 33.431744591, 14.0407622909, 62.4336607519, 5.87451869907};
test_label[1381] = '{-14.1819173741};
test_output[1381] = '{84.7579486018};
############ END DEBUG ############*/
test_input[11056:11063] = '{32'h4205fa6a, 32'hc28f4455, 32'hc149187a, 32'hc220dad0, 32'h42a9ce65, 32'h420a2ee0, 32'h42abfeed, 32'hc2035a79};
test_label[1382] = '{32'hc2035a79};
test_output[1382] = '{32'h42ee3ff2};
/*############ DEBUG ############
test_input[11056:11063] = '{33.4945432387, -71.6334581606, -12.5684753897, -40.2136834522, 84.9031132416, 34.5457767062, 85.9979007657, -32.8383519814};
test_label[1382] = '{-32.8383519814};
test_output[1382] = '{119.124892383};
############ END DEBUG ############*/
test_input[11064:11071] = '{32'hc2854fd5, 32'hc1c8177c, 32'hc137741b, 32'hc17d8d73, 32'h4118d631, 32'h41785ad5, 32'h422b61ae, 32'hbf993e00};
test_label[1383] = '{32'hbf993e00};
test_output[1383] = '{32'h42302b9e};
/*############ DEBUG ############
test_input[11064:11071] = '{-66.6559210945, -25.0114665684, -11.465845636, -15.8470332914, 9.55229270375, 15.5221753504, 42.8453888992, -1.19720464059};
test_label[1383] = '{-1.19720464059};
test_output[1383] = '{44.0425935398};
############ END DEBUG ############*/
test_input[11072:11079] = '{32'h40d7d557, 32'hc11b4846, 32'h428d8e87, 32'hc25b1f74, 32'h425049dc, 32'h41dc215f, 32'h42a2a683, 32'hc08ee94d};
test_label[1384] = '{32'hc08ee94d};
test_output[1384] = '{32'h42ab951b};
/*############ DEBUG ############
test_input[11072:11079] = '{6.74479225342, -9.70514446577, 70.7783767911, -54.7807175013, 52.0721285917, 27.5162952483, 81.3252152377, -4.46597891891};
test_label[1384] = '{-4.46597891891};
test_output[1384] = '{85.7912204326};
############ END DEBUG ############*/
test_input[11080:11087] = '{32'hc2c58e58, 32'h42865e67, 32'hc25ccbb4, 32'hc20aaa35, 32'h42958331, 32'h426a35fd, 32'h42b2eaf2, 32'h41f2baeb};
test_label[1385] = '{32'h42865e67};
test_output[1385] = '{32'h41b23229};
/*############ DEBUG ############
test_input[11080:11087] = '{-98.7780152763, 67.1843822212, -55.1989279429, -34.6662167098, 74.7562294822, 58.5527233527, 89.4588745676, 30.3412690516};
test_label[1385] = '{67.1843822212};
test_output[1385] = '{22.2744927584};
############ END DEBUG ############*/
test_input[11088:11095] = '{32'h41f28e06, 32'hc26484ad, 32'h42347be3, 32'h42819647, 32'hc1a57a26, 32'h42aa1ca2, 32'hc1dfdbe3, 32'h41be5a87};
test_label[1386] = '{32'h42347be3};
test_output[1386] = '{32'h421fbd62};
/*############ DEBUG ############
test_input[11088:11095] = '{30.3193474632, -57.129567556, 45.1209826893, 64.7935117454, -20.6846420167, 85.0559265634, -27.9823656432, 23.7942028165};
test_label[1386] = '{45.1209826893};
test_output[1386] = '{39.9349438757};
############ END DEBUG ############*/
test_input[11096:11103] = '{32'hc2a09f05, 32'hc2b4552e, 32'hc2c2d935, 32'hc016205e, 32'h424d6f11, 32'hc2b2fc94, 32'hc2746e07, 32'h42a84f03};
test_label[1387] = '{32'hc2746e07};
test_output[1387] = '{32'h43114303};
/*############ DEBUG ############
test_input[11096:11103] = '{-80.3105870001, -90.1663683071, -97.4242324097, -2.34572551662, 51.358463513, -89.4933174258, -61.1074500042, 84.1543195198};
test_label[1387] = '{-61.1074500042};
test_output[1387] = '{145.261769524};
############ END DEBUG ############*/
test_input[11104:11111] = '{32'h42b3155a, 32'h42a74cb8, 32'hc1f7babb, 32'hc1f8de5a, 32'hc2468e86, 32'h4289ded9, 32'hc2a76b23, 32'h421c8993};
test_label[1388] = '{32'h42a74cb8};
test_output[1388] = '{32'h40bca0b6};
/*############ DEBUG ############
test_input[11104:11111] = '{89.5417034969, 83.6498434701, -30.9661763672, -31.1085698239, -49.6391814665, 68.9352474829, -83.7092534986, 39.134350172};
test_label[1388] = '{83.6498434701};
test_output[1388] = '{5.89461805589};
############ END DEBUG ############*/
test_input[11112:11119] = '{32'hc18982fa, 32'h42a12020, 32'hc29ad284, 32'h42a53ca5, 32'h41244710, 32'hc0f18b08, 32'h425d987a, 32'h41f4b914};
test_label[1389] = '{32'hc0f18b08};
test_output[1389] = '{32'h42b49301};
/*############ DEBUG ############
test_input[11112:11119] = '{-17.1889533177, 80.5627425269, -77.4111629017, 82.6184467245, 10.2673492842, -7.54822150411, 55.3989030864, 30.5903710964};
test_label[1389] = '{-7.54822150411};
test_output[1389] = '{90.287116744};
############ END DEBUG ############*/
test_input[11120:11127] = '{32'hc0573ad5, 32'h41285688, 32'hc2941616, 32'hc2877445, 32'h42221c3d, 32'h418dfb73, 32'hc1048fd1, 32'h410d6686};
test_label[1390] = '{32'hc0573ad5};
test_output[1390] = '{32'h422f8feb};
/*############ DEBUG ############
test_input[11120:11127] = '{-3.36296574385, 10.5211259406, -74.0431346313, -67.7270919777, 40.5275778676, 17.7477772971, -8.28511120358, 8.83752965979};
test_label[1390] = '{-3.36296574385};
test_output[1390] = '{43.8905436116};
############ END DEBUG ############*/
test_input[11128:11135] = '{32'hc1dd6670, 32'hc29afff1, 32'h406f0c44, 32'hc2977bf3, 32'hc2b70a0c, 32'h425495c9, 32'hc22aa1f2, 32'hc2a8be1c};
test_label[1391] = '{32'hc2977bf3};
test_output[1391] = '{32'h4300e36c};
/*############ DEBUG ############
test_input[11128:11135] = '{-27.6750178341, -77.4998842475, 3.73512369941, -75.7420909722, -91.5196250542, 53.1462742518, -42.6581500098, -84.3713039343};
test_label[1391] = '{-75.7420909722};
test_output[1391] = '{128.888365224};
############ END DEBUG ############*/
test_input[11136:11143] = '{32'hc2b47a98, 32'hc262a12e, 32'hc2a7ccee, 32'hc2585be0, 32'h425ba991, 32'hc292f0a7, 32'hc1f51412, 32'h423b96a0};
test_label[1392] = '{32'hc292f0a7};
test_output[1392] = '{32'h430062cd};
/*############ DEBUG ############
test_input[11136:11143] = '{-90.2394425179, -56.6574017531, -83.9002517601, -54.0897204367, 54.9155932978, -73.4700240023, -30.6348006211, 46.8970957868};
test_label[1392] = '{-73.4700240023};
test_output[1392] = '{128.38594656};
############ END DEBUG ############*/
test_input[11144:11151] = '{32'hc12d06f0, 32'h41e6dab1, 32'hc19ec63c, 32'hc1061fea, 32'h4159a196, 32'h410ac5f3, 32'h41bd9321, 32'h42ad2243};
test_label[1393] = '{32'h42ad2243};
test_output[1393] = '{32'h80000000};
/*############ DEBUG ############
test_input[11144:11151] = '{-10.8141933698, 28.8567832758, -19.846793952, -8.38279166583, 13.6019500458, 8.6733270078, 23.6968393519, 86.5669137383};
test_label[1393] = '{86.5669137383};
test_output[1393] = '{-0.0};
############ END DEBUG ############*/
test_input[11152:11159] = '{32'hc27c4983, 32'h428e1d40, 32'h40b174e6, 32'hc2adf078, 32'h41d34b63, 32'h418f7c56, 32'hc28adc60, 32'hc24fd9d3};
test_label[1394] = '{32'hc28adc60};
test_output[1394] = '{32'h430c7cd0};
/*############ DEBUG ############
test_input[11152:11159] = '{-63.0717870731, 71.0571321848, 5.54551967553, -86.9696652571, 26.4118108678, 17.9357110827, -69.4304168892, -51.9627202865};
test_label[1394] = '{-69.4304168892};
test_output[1394] = '{140.487549074};
############ END DEBUG ############*/
test_input[11160:11167] = '{32'h41fe6517, 32'h40a48067, 32'hc22c5773, 32'hc274e594, 32'hc248a264, 32'h429d0a4f, 32'h42b8a849, 32'h42c28245};
test_label[1395] = '{32'h40a48067};
test_output[1395] = '{32'h42b83df2};
/*############ DEBUG ############
test_input[11160:11167] = '{31.7993606017, 5.14067389353, -43.0854012459, -61.2241983275, -50.1585834154, 78.5201301588, 92.3286828773, 97.2544315195};
test_label[1395] = '{5.14067389353};
test_output[1395] = '{92.120988717};
############ END DEBUG ############*/
test_input[11168:11175] = '{32'h41db49e1, 32'hc2c1f919, 32'hc2b560a0, 32'h42864d0c, 32'hc2b5726d, 32'h41f520bb, 32'hc2a2d4e7, 32'h42b7fa24};
test_label[1396] = '{32'hc2b560a0};
test_output[1396] = '{32'h4336ad62};
/*############ DEBUG ############
test_input[11168:11175] = '{27.411073504, -96.9865159492, -90.6887199541, 67.1504851182, -90.7234855333, 30.6409807773, -81.4158238905, 91.9885524316};
test_label[1396] = '{-90.6887199541};
test_output[1396] = '{182.677272386};
############ END DEBUG ############*/
test_input[11176:11183] = '{32'h420ed620, 32'hc134ce25, 32'h413de098, 32'h4163be0a, 32'hc290e5ea, 32'h413c2819, 32'h4286716d, 32'hc1784588};
test_label[1397] = '{32'h413de098};
test_output[1397] = '{32'h425d6ab3};
/*############ DEBUG ############
test_input[11176:11183] = '{35.7091046024, -11.3003279816, 11.8673325897, 14.2338966008, -72.4490478919, 11.7597898445, 67.2215319281, -15.5169751609};
test_label[1397] = '{11.8673325897};
test_output[1397] = '{55.3541993384};
############ END DEBUG ############*/
test_input[11184:11191] = '{32'hc166098a, 32'hc0570b45, 32'h42949cc1, 32'h42385f60, 32'hc17cc286, 32'h42bbcef1, 32'hc258c448, 32'hc2bb03bf};
test_label[1398] = '{32'h42949cc1};
test_output[1398] = '{32'h419cc8c2};
/*############ DEBUG ############
test_input[11184:11191] = '{-14.3773285395, -3.36006279581, 74.3061582174, 46.0931411825, -15.7974908044, 93.9041838732, -54.1916801563, -93.507314872};
test_label[1398] = '{74.3061582174};
test_output[1398] = '{19.5980256589};
############ END DEBUG ############*/
test_input[11192:11199] = '{32'h424c1be7, 32'h425083ae, 32'hc2b711d7, 32'h42a56996, 32'hc1def589, 32'hc1844a97, 32'h41cdc395, 32'h42938d2f};
test_label[1399] = '{32'hc2b711d7};
test_output[1399] = '{32'h432e3dbf};
/*############ DEBUG ############
test_input[11192:11199] = '{51.0272494505, 52.128595075, -91.5348419438, 82.7062187292, -27.8698899941, -16.5364213925, 25.7204999633, 73.7757464798};
test_label[1399] = '{-91.5348419438};
test_output[1399] = '{174.24119296};
############ END DEBUG ############*/
test_input[11200:11207] = '{32'h42c222b9, 32'hc15e4cdf, 32'hc24d3c64, 32'hc2c3ab86, 32'hc2bb1ef3, 32'h422506bd, 32'hc2acf624, 32'hc081ae7a};
test_label[1400] = '{32'h42c222b9};
test_output[1400] = '{32'h80000000};
/*############ DEBUG ############
test_input[11200:11207] = '{97.0678190766, -13.8937670572, -51.3089765455, -97.8350036208, -93.5604445487, 41.2565810422, -86.4807430691, -4.05254824872};
test_label[1400] = '{97.0678190766};
test_output[1400] = '{-0.0};
############ END DEBUG ############*/
test_input[11208:11215] = '{32'h418b1a91, 32'h424e1b58, 32'h42277285, 32'h4284b726, 32'hc199ab81, 32'h41a8d771, 32'hc2931074, 32'hc2620cf2};
test_label[1401] = '{32'h4284b726};
test_output[1401] = '{32'h34c27a68};
/*############ DEBUG ############
test_input[11208:11215] = '{17.387972021, 51.5267015438, 41.8618337039, 66.35771322, -19.2087415449, 21.1051967154, -73.5321363852, -56.5126409137};
test_label[1401] = '{66.35771322};
test_output[1401] = '{3.62243795178e-07};
############ END DEBUG ############*/
test_input[11216:11223] = '{32'h422549be, 32'hc2446731, 32'hc17f1079, 32'hc212a5e2, 32'h429f28cb, 32'h42c04ae4, 32'h42601144, 32'hc2822f0a};
test_label[1402] = '{32'h422549be};
test_output[1402] = '{32'h425b4c0a};
/*############ DEBUG ############
test_input[11216:11223] = '{41.3220128908, -49.1007730116, -15.9415212087, -36.6619934769, 79.5796736024, 96.146269573, 56.0168623312, -65.0918733989};
test_label[1402] = '{41.3220128908};
test_output[1402] = '{54.8242567461};
############ END DEBUG ############*/
test_input[11224:11231] = '{32'h4206eda0, 32'h428693d3, 32'h421ffd41, 32'hc2802f3f, 32'h4295c055, 32'h411fd76a, 32'hc2a4ef82, 32'hc1fdfefd};
test_label[1403] = '{32'h411fd76a};
test_output[1403] = '{32'h4281c5aa};
/*############ DEBUG ############
test_input[11224:11231] = '{33.7320559815, 67.288716499, 39.9973188652, -64.0922781695, 74.8756470979, 9.99009099461, -82.4677893943, -31.7495052836};
test_label[1403] = '{9.99009099461};
test_output[1403] = '{64.8860630098};
############ END DEBUG ############*/
test_input[11232:11239] = '{32'h42c7951a, 32'hc2adb311, 32'h42bd1452, 32'h4294453e, 32'h4220322d, 32'h4206326f, 32'h3f65aee3, 32'hc23275f6};
test_label[1404] = '{32'h42bd1452};
test_output[1404] = '{32'h40a83754};
/*############ DEBUG ############
test_input[11232:11239] = '{99.7912143712, -86.8497379967, 94.5396861098, 74.1352400375, 40.0490006388, 33.5492526425, 0.897199790512, -44.6151970424};
test_label[1404] = '{94.5396861098};
test_output[1404] = '{5.25675408791};
############ END DEBUG ############*/
test_input[11240:11247] = '{32'hc2b007af, 32'h42702035, 32'h41748812, 32'hc1200a2a, 32'h41aad735, 32'h42687f3d, 32'h41b690f1, 32'h42a983f8};
test_label[1405] = '{32'h42a983f8};
test_output[1405] = '{32'h2db87840};
/*############ DEBUG ############
test_input[11240:11247] = '{-88.0150060127, 60.0314527244, 15.2832201167, -10.0024814281, 21.3550810301, 58.1242554301, 22.8207718903, 84.7577484823};
test_label[1405] = '{84.7577484823};
test_output[1405] = '{2.09717798685e-11};
############ END DEBUG ############*/
test_input[11248:11255] = '{32'h428ecf1c, 32'hc1e595b0, 32'hc149a878, 32'hc2c471d7, 32'h428849c8, 32'hc2aa7d5c, 32'hc29ed413, 32'hc265f707};
test_label[1406] = '{32'hc2aa7d5c};
test_output[1406] = '{32'h431cafe0};
/*############ DEBUG ############
test_input[11248:11255] = '{71.4045077148, -28.6980896386, -12.6036299788, -98.2223410724, 68.1441064376, -85.2448442325, -79.4142105506, -57.4912367309};
test_label[1406] = '{-85.2448442325};
test_output[1406] = '{156.687007009};
############ END DEBUG ############*/
test_input[11256:11263] = '{32'hc1d136ec, 32'hc1f7abca, 32'h4062efad, 32'hc2938f5d, 32'h410783ea, 32'hc2c68475, 32'hc2bf8458, 32'hc0f51fc3};
test_label[1407] = '{32'hc0f51fc3};
test_output[1407] = '{32'h418118bc};
/*############ DEBUG ############
test_input[11256:11263] = '{-26.1518164229, -30.9588820004, 3.54587863093, -73.7800053317, 8.46970547244, -99.2587032259, -95.7584833467, -7.66012725984};
test_label[1407] = '{-7.66012725984};
test_output[1407] = '{16.1370777739};
############ END DEBUG ############*/
test_input[11264:11271] = '{32'h4285d727, 32'h424fd122, 32'h408ec381, 32'hc1863a25, 32'hc2bc7b7e, 32'h3f9ede90, 32'h421e9b9d, 32'hc1d344a6};
test_label[1408] = '{32'h3f9ede90};
test_output[1408] = '{32'h42835bad};
/*############ DEBUG ############
test_input[11264:11271] = '{66.9202226013, 51.9542328282, 4.46136516122, -16.7783901219, -94.2411954949, 1.24116703927, 39.6519652224, -26.4085192198};
test_label[1408] = '{1.24116703927};
test_output[1408] = '{65.6790558785};
############ END DEBUG ############*/
test_input[11272:11279] = '{32'h41e1afe9, 32'h4235cd32, 32'h42a84963, 32'h4080c593, 32'hc269276a, 32'hc2500e28, 32'hc2a7ddb3, 32'hc18f291f};
test_label[1409] = '{32'h4080c593};
test_output[1409] = '{32'h42a03d0a};
/*############ DEBUG ############
test_input[11272:11279] = '{28.2108929659, 45.4503864172, 84.1433354945, 4.02411785406, -58.2884910696, -52.0138239205, -83.9330072753, -17.8950793184};
test_label[1409] = '{4.02411785406};
test_output[1409] = '{80.1192176404};
############ END DEBUG ############*/
test_input[11280:11287] = '{32'h42aa8d14, 32'h417b66b6, 32'h422e5009, 32'hc1af5702, 32'hc2bca4f8, 32'h424a8508, 32'h40b5b4cf, 32'hc2a4c96f};
test_label[1410] = '{32'h424a8508};
test_output[1410] = '{32'h420a9520};
/*############ DEBUG ############
test_input[11280:11287] = '{85.2755441125, 15.7125754384, 43.5781599757, -21.9174837834, -94.322203232, 50.6299146367, 5.67832126357, -82.3934237946};
test_label[1410] = '{50.6299146367};
test_output[1410] = '{34.6456294758};
############ END DEBUG ############*/
test_input[11288:11295] = '{32'h41a0b4ee, 32'h413dca35, 32'h419d7990, 32'h42af4aa8, 32'hc20d8dd4, 32'h4267421c, 32'hc2be443e, 32'h42b56886};
test_label[1411] = '{32'hc2be443e};
test_output[1411] = '{32'h4339e222};
/*############ DEBUG ############
test_input[11288:11295] = '{20.088344282, 11.8618665511, 19.6843564983, 87.645811523, -35.3885037499, 57.8145599902, -95.1332823147, 90.7041473169};
test_label[1411] = '{-95.1332823147};
test_output[1411] = '{185.88332589};
############ END DEBUG ############*/
test_input[11296:11303] = '{32'h429609ef, 32'hc0ef62d2, 32'hc2393d82, 32'hc296c6cf, 32'h42405b9f, 32'h417ffa0f, 32'h428b613b, 32'h42769bfb};
test_label[1412] = '{32'h42769bfb};
test_output[1412] = '{32'h4155f35d};
/*############ DEBUG ############
test_input[11296:11303] = '{75.0194032108, -7.48081315475, -46.3100674488, -75.3883003276, 48.0894729491, 15.9985498537, 69.6899069807, 61.6523246617};
test_label[1412] = '{61.6523246617};
test_output[1412] = '{13.3719149117};
############ END DEBUG ############*/
test_input[11304:11311] = '{32'hc29fb2cb, 32'h425302c2, 32'h421e96b8, 32'hc21797b7, 32'h412127b1, 32'hc2239232, 32'hc20812f8, 32'hc26a0fe2};
test_label[1413] = '{32'h425302c2};
test_output[1413] = '{32'h36087fde};
/*############ DEBUG ############
test_input[11304:11311] = '{-79.8492083338, 52.7526929544, 39.6471881158, -37.8981604354, 10.0721900836, -40.8927693426, -34.0185238427, -58.5155095137};
test_label[1413] = '{52.7526929544};
test_output[1413] = '{2.03400082323e-06};
############ END DEBUG ############*/
test_input[11312:11319] = '{32'hc13afe8d, 32'h405ec60e, 32'h4255054b, 32'hc29ec026, 32'hc26cce33, 32'h4258e6fe, 32'h428e3610, 32'h4265167a};
test_label[1414] = '{32'hc29ec026};
test_output[1414] = '{32'h43167b1b};
/*############ DEBUG ############
test_input[11312:11319] = '{-11.6871463454, 3.48083820501, 53.2551674426, -79.3752899056, -59.2013646855, 54.2255781282, 71.1055933651, 57.2719514007};
test_label[1414] = '{-79.3752899056};
test_output[1414] = '{150.480884317};
############ END DEBUG ############*/
test_input[11320:11327] = '{32'hc21c96ae, 32'hc1f10194, 32'h42ab973d, 32'h41b43fc4, 32'h42ada839, 32'hc261ae1e, 32'hc25b8290, 32'hc1194b77};
test_label[1415] = '{32'hc261ae1e};
test_output[1415] = '{32'h430f8d94};
/*############ DEBUG ############
test_input[11320:11327] = '{-39.1471475437, -30.1257698268, 85.79538583, 22.5311352969, 86.8285592711, -56.4200364064, -54.8775025639, -9.58092376542};
test_label[1415] = '{-56.4200364064};
test_output[1415] = '{143.553043282};
############ END DEBUG ############*/
test_input[11328:11335] = '{32'h42a5d083, 32'hbf8fc6c0, 32'hc2b5e4d3, 32'hc1b016af, 32'h40f79dc7, 32'h42413a02, 32'hc0d3e495, 32'hc2467839};
test_label[1416] = '{32'hc2b5e4d3};
test_output[1416] = '{32'h432ddaab};
/*############ DEBUG ############
test_input[11328:11335] = '{82.9072510061, -1.12325290459, -90.9469228892, -22.0110750883, 7.73800985927, 48.3066492215, -6.62165319076, -49.6174058081};
test_label[1416] = '{-90.9469228892};
test_output[1416] = '{173.854173895};
############ END DEBUG ############*/
test_input[11336:11343] = '{32'hc14c9519, 32'hc294b47a, 32'hc21d3182, 32'h42892035, 32'h429d3e83, 32'hc25b9418, 32'hc1201a0a, 32'h426bfa77};
test_label[1417] = '{32'hc14c9519};
test_output[1417] = '{32'h42b6d12c};
/*############ DEBUG ############
test_input[11336:11343] = '{-12.786400455, -74.3524922694, -39.2983457707, 68.5629038913, 78.6220917963, -54.8946242755, -10.0063575864, 58.9945961594};
test_label[1417] = '{-12.786400455};
test_output[1417] = '{91.4085350442};
############ END DEBUG ############*/
test_input[11344:11351] = '{32'h41bdd565, 32'hc20684be, 32'hbf8f9842, 32'hc2579920, 32'hc2aa9c92, 32'h415fa006, 32'hc1408ae0, 32'h4258b7a7};
test_label[1418] = '{32'h415fa006};
test_output[1418] = '{32'h4220cfa6};
/*############ DEBUG ############
test_input[11344:11351] = '{23.7291963439, -33.6296310972, -1.12183407084, -53.8995350039, -85.3058013338, 13.9765678034, -12.0339051089, 54.1793482937};
test_label[1418] = '{13.9765678034};
test_output[1418] = '{40.2027804903};
############ END DEBUG ############*/
test_input[11352:11359] = '{32'hc294ac15, 32'hc26df676, 32'h42723c6b, 32'h419b488d, 32'h429caa33, 32'hc2c54810, 32'hc1b0a99c, 32'hc1b3c9df};
test_label[1419] = '{32'hc294ac15};
test_output[1419] = '{32'h4318ab24};
/*############ DEBUG ############
test_input[11352:11359] = '{-74.3360951292, -59.4906842948, 60.5590023116, 19.4104244598, 78.3324221003, -98.6407464846, -22.0828168088, -22.4735704901};
test_label[1419] = '{-74.3360951292};
test_output[1419] = '{152.668517249};
############ END DEBUG ############*/
test_input[11360:11367] = '{32'hc2bf12fe, 32'hc20c2c76, 32'h4222927f, 32'h42a1cd36, 32'hc2823a0c, 32'hc29182cb, 32'hc2b679fe, 32'hc1647d05};
test_label[1420] = '{32'hc20c2c76};
test_output[1420] = '{32'h42e7e371};
/*############ DEBUG ############
test_input[11360:11367] = '{-95.5370940246, -35.0434175739, 40.6430610331, 80.9008057998, -65.1133764871, -72.755457262, -91.238266555, -14.2805223303};
test_label[1420] = '{-35.0434175739};
test_output[1420] = '{115.944223374};
############ END DEBUG ############*/
test_input[11368:11375] = '{32'h42630ad7, 32'hc2ac96c4, 32'h429b6702, 32'hc20a728f, 32'hc20ef58e, 32'hc2b8d386, 32'hc2ad10ec, 32'h41f1967f};
test_label[1421] = '{32'hc20ef58e};
test_output[1421] = '{32'h42e2e1c9};
/*############ DEBUG ############
test_input[11368:11375] = '{56.7605840042, -86.2944676401, 77.7011884952, -34.6118749547, -35.7398000938, -92.4131320344, -86.5330542475, 30.1984837493};
test_label[1421] = '{-35.7398000938};
test_output[1421] = '{113.44098859};
############ END DEBUG ############*/
test_input[11376:11383] = '{32'h40f48b80, 32'h418dddfc, 32'h41acf607, 32'hc2a6a6b3, 32'h42233dcc, 32'hc2687adc, 32'hc2c66b57, 32'h429f2cba};
test_label[1422] = '{32'h418dddfc};
test_output[1422] = '{32'h42776a77};
/*############ DEBUG ############
test_input[11376:11383] = '{7.64202888341, 17.7333905006, 21.620130691, -83.3255881767, 40.8103472068, -58.1199787043, -99.2096472712, 79.5873582602};
test_label[1422] = '{17.7333905006};
test_output[1422] = '{61.8539677596};
############ END DEBUG ############*/
test_input[11384:11391] = '{32'h426bfd33, 32'hc1b9227a, 32'hc09a8af9, 32'h42723ab0, 32'h428dfe7c, 32'hc28afd46, 32'hbdac928f, 32'h4296d1c3};
test_label[1423] = '{32'h428dfe7c};
test_output[1423] = '{32'h408d971e};
/*############ DEBUG ############
test_input[11384:11391] = '{58.9972657375, -23.1418349529, -4.8294643107, 60.5573104478, 70.9970423499, -69.4946746918, -0.0842639102666, 75.4096888463};
test_label[1423] = '{70.9970423499};
test_output[1423] = '{4.42469707693};
############ END DEBUG ############*/
test_input[11392:11399] = '{32'hc292f8cb, 32'h42b854ef, 32'h41d1c15e, 32'h42c0921b, 32'hc298f874, 32'h423e38df, 32'h429b1509, 32'h4272f494};
test_label[1424] = '{32'h429b1509};
test_output[1424] = '{32'h4196154f};
/*############ DEBUG ############
test_input[11392:11399] = '{-73.4859214122, 92.1658889835, 26.2194183212, 96.2853638251, -76.4852625468, 47.5555363694, 77.5410821999, 60.7388451597};
test_label[1424] = '{77.5410821999};
test_output[1424] = '{18.760404013};
############ END DEBUG ############*/
test_input[11400:11407] = '{32'hc15840db, 32'hc2bd7680, 32'hc004e931, 32'h42b56cf0, 32'hc177d075, 32'h3fcdaa67, 32'h41b74457, 32'hc1b09ab1};
test_label[1425] = '{32'hc004e931};
test_output[1425] = '{32'h42b9943a};
/*############ DEBUG ############
test_input[11400:11407] = '{-13.5158338555, -94.7314475011, -2.07673283025, 90.7127715602, -15.4883928369, 1.60676274741, 22.9083691641, -22.0755319777};
test_label[1425] = '{-2.07673283025};
test_output[1425] = '{92.7895043905};
############ END DEBUG ############*/
test_input[11408:11415] = '{32'hc29c458f, 32'hc2a646fc, 32'hc2c42984, 32'hc21d342d, 32'hc2bfbb9c, 32'h42a53252, 32'h428a5324, 32'h42736816};
test_label[1426] = '{32'hc21d342d};
test_output[1426] = '{32'h42f3cc68};
/*############ DEBUG ############
test_input[11408:11415] = '{-78.135853718, -83.1386411993, -98.0810888082, -39.3009513154, -95.8664271291, 82.5982817691, 69.1623810564, 60.8516466746};
test_label[1426] = '{-39.3009513154};
test_output[1426] = '{121.899234547};
############ END DEBUG ############*/
test_input[11416:11423] = '{32'hc23fabb3, 32'hc2b8d693, 32'h421115bc, 32'h42b6c169, 32'h4153d077, 32'hc29a51d8, 32'hc2b603b1, 32'hc24678d8};
test_label[1427] = '{32'hc2b603b1};
test_output[1427] = '{32'h4336628d};
/*############ DEBUG ############
test_input[11416:11423] = '{-47.9176743323, -92.4190914772, 36.2712247526, 91.3777522654, 13.2383949355, -77.1598519232, -91.0072090402, -49.618012708};
test_label[1427] = '{-91.0072090402};
test_output[1427] = '{182.384961306};
############ END DEBUG ############*/
test_input[11424:11431] = '{32'hc0ba939f, 32'h427740ba, 32'hc2507d5c, 32'hbf507bcd, 32'h425ab1b4, 32'h42a9bcaa, 32'hc20541d7, 32'hc21c38a7};
test_label[1428] = '{32'hc21c38a7};
test_output[1428] = '{32'h42f7d8fe};
/*############ DEBUG ############
test_input[11424:11431] = '{-5.83052019459, 61.813210323, -52.1224198032, -0.81438903443, 54.6735391851, 84.8684855656, -33.3142957303, -39.0553242867};
test_label[1428] = '{-39.0553242867};
test_output[1428] = '{123.923809852};
############ END DEBUG ############*/
test_input[11432:11439] = '{32'h4205365c, 32'hc2ba31a8, 32'h4269934c, 32'h423d773d, 32'hc269f781, 32'hc1a679ce, 32'hc1e9e55d, 32'h419e1f0b};
test_label[1429] = '{32'hc2ba31a8};
test_output[1429] = '{32'h43177da8};
/*############ DEBUG ############
test_input[11432:11439] = '{33.3030836957, -93.096987932, 58.3938461641, 47.3664429255, -58.4917028784, -20.8094750249, -29.236994356, 19.7651583047};
test_label[1429] = '{-93.096987932};
test_output[1429] = '{151.490850346};
############ END DEBUG ############*/
test_input[11440:11447] = '{32'hc25aa316, 32'hc27bf000, 32'h41cb375b, 32'h410911ae, 32'h416da791, 32'h42819c39, 32'h4288cbcf, 32'hc13e1a11};
test_label[1430] = '{32'h416da791};
test_output[1430] = '{32'h42564985};
/*############ DEBUG ############
test_input[11440:11447] = '{-54.6592652211, -62.9843741425, 25.4020293827, 8.56681589626, 14.8534100171, 64.8051239402, 68.3980625371, -11.8813640026};
test_label[1430] = '{14.8534100171};
test_output[1430] = '{53.5717980721};
############ END DEBUG ############*/
test_input[11448:11455] = '{32'h42141c27, 32'h4261e9b2, 32'hc215cb2f, 32'hc2557bb2, 32'hc01997a7, 32'h429b8a4b, 32'h42595638, 32'hc1e95d5d};
test_label[1431] = '{32'h42595638};
test_output[1431] = '{32'h41bb7cbb};
/*############ DEBUG ############
test_input[11448:11455] = '{37.0274923722, 56.4782196005, -37.4484216207, -53.3707953474, -2.39988107555, 77.7701013259, 54.3341985133, -29.1705883889};
test_label[1431] = '{54.3341985133};
test_output[1431] = '{23.4359028132};
############ END DEBUG ############*/
test_input[11456:11463] = '{32'hc21cc2b6, 32'hc1957887, 32'h4175c306, 32'h41e0918c, 32'hc00c7969, 32'hc2acd2a4, 32'h419bf170, 32'hc2906692};
test_label[1432] = '{32'hc00c7969};
test_output[1432] = '{32'h41f2211d};
/*############ DEBUG ############
test_input[11456:11463] = '{-39.1901468618, -18.6838509248, 15.3601135691, 28.0710668699, -2.19491027348, -86.4114052918, 19.4928890237, -72.2003363683};
test_label[1432] = '{-2.19491027348};
test_output[1432] = '{30.2661683105};
############ END DEBUG ############*/
test_input[11464:11471] = '{32'h3fac14ae, 32'hc2b934bd, 32'h42961a21, 32'hc1df9d86, 32'hc23075ad, 32'h4293235b, 32'hbf76fd77, 32'h424e0c28};
test_label[1433] = '{32'hc1df9d86};
test_output[1433] = '{32'h42ce6a54};
/*############ DEBUG ############
test_input[11464:11471] = '{1.3443810704, -92.6030062203, 75.0510312792, -27.951914853, -44.1149164268, 73.5690524317, -0.964805062714, 51.5118696197};
test_label[1433] = '{-27.951914853};
test_output[1433] = '{103.207671239};
############ END DEBUG ############*/
test_input[11472:11479] = '{32'hc01c3737, 32'hc1d6c6e4, 32'hc2b7e7ff, 32'h422b7d78, 32'hc2a16921, 32'h41275d93, 32'h4282a179, 32'hc1f16915};
test_label[1434] = '{32'h422b7d78};
test_output[1434] = '{32'h41b38af3};
/*############ DEBUG ############
test_input[11472:11479] = '{-2.44086997721, -26.8471149842, -91.9531135999, 42.8725285474, -80.7053295109, 10.460345686, 65.3153745604, -30.1763094087};
test_label[1434] = '{42.8725285474};
test_output[1434] = '{22.4428460132};
############ END DEBUG ############*/
test_input[11480:11487] = '{32'h423917f3, 32'h428c0030, 32'hc2076e6b, 32'hc284fc0a, 32'hc2c0e787, 32'hc2a9e747, 32'hc2860fa3, 32'hc2b6856b};
test_label[1435] = '{32'h423917f3};
test_output[1435] = '{32'h41bdd0d9};
/*############ DEBUG ############
test_input[11480:11487] = '{46.2733888615, 70.0003646804, -33.8578312595, -66.4922638343, -96.4522015299, -84.9517165469, -67.0305439298, -91.2605808527};
test_label[1435] = '{46.2733888615};
test_output[1435] = '{23.726975819};
############ END DEBUG ############*/
test_input[11488:11495] = '{32'h420ded02, 32'h42983004, 32'h415f2fd7, 32'h4234d3fc, 32'hc26571c1, 32'hc2a81f98, 32'hbdd007db, 32'hc1132b12};
test_label[1436] = '{32'h415f2fd7};
test_output[1436] = '{32'h42789411};
/*############ DEBUG ############
test_input[11488:11495] = '{35.4814516128, 76.0937769465, 13.9491793305, 45.2070173923, -57.361086109, -84.0617096193, -0.101577481058, -9.19801485435};
test_label[1436] = '{13.9491793305};
test_output[1436] = '{62.144597616};
############ END DEBUG ############*/
test_input[11496:11503] = '{32'hc0790257, 32'hc2041793, 32'h41f4b6b0, 32'h42c7d96d, 32'hc24410b2, 32'h40ca7e1e, 32'h423b605d, 32'h4244d230};
test_label[1437] = '{32'h42c7d96d};
test_output[1437] = '{32'h80000000};
/*############ DEBUG ############
test_input[11496:11503] = '{-3.89076779892, -33.0230227323, 30.5892036576, 99.9246604227, -49.0163057322, 6.32789502969, 46.8441052217, 49.2052620684};
test_label[1437] = '{99.9246604227};
test_output[1437] = '{-0.0};
############ END DEBUG ############*/
test_input[11504:11511] = '{32'h41ea369d, 32'h42b79c24, 32'h42b1245c, 32'hc1492285, 32'hc2c6effe, 32'h4170ba57, 32'h427dc80b, 32'hc20060f3};
test_label[1438] = '{32'h427dc80b};
test_output[1438] = '{32'h41e32f9e};
/*############ DEBUG ############
test_input[11504:11511] = '{29.2766658065, 91.8049596424, 88.5710128498, -12.5709274345, -99.4687343673, 15.0454934364, 63.4453550474, -32.0946776054};
test_label[1438] = '{63.4453550474};
test_output[1438] = '{28.3982498361};
############ END DEBUG ############*/
test_input[11512:11519] = '{32'h3fc15b4f, 32'h41d8976a, 32'hc190ea6c, 32'hc193ebc5, 32'h428809c2, 32'hc1ae76a5, 32'h42b15e30, 32'hc131810f};
test_label[1439] = '{32'hc190ea6c};
test_output[1439] = '{32'h42d598cc};
/*############ DEBUG ############
test_input[11512:11519] = '{1.51059898524, 27.0739319343, -18.114464357, -18.4901211195, 68.0190573368, -21.8079319712, 88.683963487, -11.0940089017};
test_label[1439] = '{-18.114464357};
test_output[1439] = '{106.798427845};
############ END DEBUG ############*/
test_input[11520:11527] = '{32'hc273bf13, 32'hc225fdc6, 32'h408187b8, 32'h424b6ca3, 32'h42a40c42, 32'h42bdd6c3, 32'h40c16f06, 32'h3ff7dfa1};
test_label[1440] = '{32'h42a40c42};
test_output[1440] = '{32'h414e540a};
/*############ DEBUG ############
test_input[11520:11527] = '{-60.9365967803, -41.4978240623, 4.04781733735, 50.8560915223, 82.0239388648, 94.9194538176, 6.04480264534, 1.93651216246};
test_label[1440] = '{82.0239388648};
test_output[1440] = '{12.8955174621};
############ END DEBUG ############*/
test_input[11528:11535] = '{32'h40f44580, 32'hc2a0c9df, 32'h425d21f6, 32'hc2b71771, 32'hc2a50a6c, 32'hc271a235, 32'hc2b7680e, 32'hc2a9151b};
test_label[1441] = '{32'hc2a0c9df};
test_output[1441] = '{32'h4307ad6d};
/*############ DEBUG ############
test_input[11528:11535] = '{7.63348388879, -80.3942775505, 55.2831635193, -91.5457855598, -82.5203517527, -60.4084045361, -91.7032297462, -84.5412242974};
test_label[1441] = '{-80.3942775505};
test_output[1441] = '{135.67744107};
############ END DEBUG ############*/
test_input[11536:11543] = '{32'h42ac1440, 32'hc2150c6e, 32'hc1fd18f7, 32'hbfa40067, 32'hc0e940b4, 32'h4263d166, 32'hc1e3327e, 32'hc20b736c};
test_label[1442] = '{32'hc1fd18f7};
test_output[1442] = '{32'h42eb5a7d};
/*############ DEBUG ############
test_input[11536:11543] = '{86.0395475897, -37.2621372599, -31.6371904303, -1.28126225856, -7.28914853995, 56.9544910846, -28.399654354, -34.8627160287};
test_label[1442] = '{-31.6371904303};
test_output[1442] = '{117.67673802};
############ END DEBUG ############*/
test_input[11544:11551] = '{32'hc195b06f, 32'h42c36594, 32'hc1c8bad1, 32'h4185e246, 32'h41038158, 32'h3fe57fc1, 32'h42747493, 32'h4082961c};
test_label[1443] = '{32'h4185e246};
test_output[1443] = '{32'h42a1ed02};
/*############ DEBUG ############
test_input[11544:11551] = '{-18.7111487244, 97.698393739, -25.0912194923, 16.7354853206, 8.21907766483, 1.79296125669, 61.1138408724, 4.08082410156};
test_label[1443] = '{16.7354853206};
test_output[1443] = '{80.9629084185};
############ END DEBUG ############*/
test_input[11552:11559] = '{32'h428fb466, 32'hc27c1063, 32'hc2ac1718, 32'h42c0725d, 32'h42963d2e, 32'h429d8456, 32'h42b150f3, 32'h418a9fd9};
test_label[1444] = '{32'h42963d2e};
test_output[1444] = '{32'h41a8d5cb};
/*############ DEBUG ############
test_input[11552:11559] = '{71.8523386344, -63.0160016541, -86.0451068143, 96.2233664385, 75.1194937285, 78.7584701845, 88.658100696, 17.3280512551};
test_label[1444] = '{75.1194937285};
test_output[1444] = '{21.1043907421};
############ END DEBUG ############*/
test_input[11560:11567] = '{32'hc24fc252, 32'h425e6f0c, 32'hc2a187d4, 32'hc208baf1, 32'hc10bcde5, 32'h428d4447, 32'hc1c36fda, 32'hc2904b9e};
test_label[1445] = '{32'hc10bcde5};
test_output[1445] = '{32'h429ebe04};
/*############ DEBUG ############
test_input[11560:11567] = '{-51.9397642019, 55.6084434144, -80.7652887219, -34.1825611195, -8.73776741685, 70.6333561566, -24.429615259, -72.1476876451};
test_label[1445] = '{-8.73776741685};
test_output[1445] = '{79.3711238719};
############ END DEBUG ############*/
test_input[11568:11575] = '{32'hc2333fc0, 32'h429c80fb, 32'h42086c05, 32'h428c503f, 32'h3ffa3809, 32'h4234ddc4, 32'hc235c90a, 32'hc29bada8};
test_label[1446] = '{32'h42086c05};
test_output[1446] = '{32'h42309641};
/*############ DEBUG ############
test_input[11568:11575] = '{-44.8122564843, 78.2519167874, 34.1054885252, 70.1567276565, 1.95483499863, 45.2165669835, -45.4463286065, -77.8391686534};
test_label[1446] = '{34.1054885252};
test_output[1446] = '{44.1467332187};
############ END DEBUG ############*/
test_input[11576:11583] = '{32'hc1fd281e, 32'hc28eba5f, 32'h42519e45, 32'hc2abd34c, 32'h41ce236a, 32'h42a69df1, 32'h3fd3e5af, 32'hc07b7cd5};
test_label[1447] = '{32'h42519e45};
test_output[1447] = '{32'h41f73b3c};
/*############ DEBUG ############
test_input[11576:11583] = '{-31.6445879309, -71.3640028511, 52.4045588796, -85.9126868932, 25.7672918527, 83.3084824612, 1.65544694369, -3.92949412111};
test_label[1447] = '{52.4045588796};
test_output[1447] = '{30.9039235817};
############ END DEBUG ############*/
test_input[11584:11591] = '{32'hc25b3d0f, 32'hc1b53984, 32'h41bfda5e, 32'h4246a754, 32'h4246fdb5, 32'hc2799a0d, 32'hc168bcf1, 32'hc28c7cc9};
test_label[1448] = '{32'hc25b3d0f};
test_output[1448] = '{32'h42d26b23};
/*############ DEBUG ############
test_input[11584:11591] = '{-54.8096291584, -22.6530842601, 23.9816237853, 49.6634061784, 49.7477596092, -62.4004420799, -14.5461283635, -70.2437184594};
test_label[1448] = '{-54.8096291584};
test_output[1448] = '{105.209248407};
############ END DEBUG ############*/
test_input[11592:11599] = '{32'h4162a089, 32'hc1ba91c7, 32'h421cb350, 32'h3ef1ff82, 32'hc1d0c7ca, 32'h4207939e, 32'hc22ea867, 32'hc06da865};
test_label[1449] = '{32'hc22ea867};
test_output[1449] = '{32'h42a5b075};
/*############ DEBUG ############
test_input[11592:11599] = '{14.1641930833, -23.321181287, 39.1751094165, 0.472652487745, -26.0975540857, 33.8941577527, -43.664454733, -3.71340309363};
test_label[1449] = '{-43.664454733};
test_output[1449] = '{82.8446388383};
############ END DEBUG ############*/
test_input[11600:11607] = '{32'hc27f2579, 32'h422eea52, 32'hc2a98c67, 32'hc2971d31, 32'h4022d7fa, 32'h4290421e, 32'h42c0bbb8, 32'h42c4aa3c};
test_label[1450] = '{32'hc2971d31};
test_output[1450] = '{32'h432e0544};
/*############ DEBUG ############
test_input[11600:11607] = '{-63.7865960079, 43.728827506, -84.7742226403, -75.5570166882, 2.54443206145, 72.129136582, 96.3666372864, 98.3324884359};
test_label[1450] = '{-75.5570166882};
test_output[1450] = '{174.02056553};
############ END DEBUG ############*/
test_input[11608:11615] = '{32'h41b1f779, 32'h41048ae6, 32'h41c48f68, 32'hc195321e, 32'h4243a61d, 32'hc2a44722, 32'hc28a1994, 32'h410a2d3e};
test_label[1451] = '{32'hc2a44722};
test_output[1451] = '{32'h43030d18};
/*############ DEBUG ############
test_input[11608:11615] = '{22.2458362466, 8.28391110237, 24.5700232264, -18.6494712994, 48.9122205311, -82.138929298, -69.0499609133, 8.6360452667};
test_label[1451] = '{-82.138929298};
test_output[1451] = '{131.051149829};
############ END DEBUG ############*/
test_input[11616:11623] = '{32'h42a1901f, 32'hc08ab850, 32'h41cebe3d, 32'hc295a329, 32'h4256d91a, 32'h4209d0d9, 32'h415cb201, 32'h42887c0d};
test_label[1452] = '{32'hc295a329};
test_output[1452] = '{32'h431b99a5};
/*############ DEBUG ############
test_input[11616:11623] = '{80.7814882005, -4.33499903336, 25.8428891643, -74.8186752274, 53.7120139237, 34.4539517332, 13.7934584407, 68.2422895969};
test_label[1452] = '{-74.8186752274};
test_output[1452] = '{155.600167011};
############ END DEBUG ############*/
test_input[11624:11631] = '{32'h42aa72ab, 32'h42227e50, 32'hc1b60862, 32'hc157a4d4, 32'h42a1ba31, 32'h421f30a5, 32'h423306ff, 32'h42aa461a};
test_label[1453] = '{32'h42aa72ab};
test_output[1453] = '{32'h3f283f49};
/*############ DEBUG ############
test_input[11624:11631] = '{85.2239606205, 40.6233510881, -22.7540933977, -13.4777410167, 80.8636527977, 39.7975063306, 44.7568306698, 85.1369182381};
test_label[1453] = '{85.2239606205};
test_output[1453] = '{0.657215656185};
############ END DEBUG ############*/
test_input[11632:11639] = '{32'hc2b35001, 32'h42c5d392, 32'hc1851e48, 32'hc1fdf6a5, 32'hc21225ab, 32'h42bd831b, 32'hc29cab81, 32'h42733b40};
test_label[1454] = '{32'h42733b40};
test_output[1454] = '{32'h42187bca};
/*############ DEBUG ############
test_input[11632:11639] = '{-89.6562591343, 98.9132205172, -16.6397864075, -31.745431961, -36.5367835829, 94.7560668901, -78.3349676965, 60.8078625256};
test_label[1454] = '{60.8078625256};
test_output[1454] = '{38.1208888078};
############ END DEBUG ############*/
test_input[11640:11647] = '{32'hc2a28267, 32'hc254582d, 32'hc1c03764, 32'hc084d1af, 32'hc07b1e8c, 32'hc26d766b, 32'h419dd9f2, 32'hc2c0ef0a};
test_label[1455] = '{32'h419dd9f2};
test_output[1455] = '{32'h2ed29c80};
/*############ DEBUG ############
test_input[11640:11647] = '{-81.2546945039, -53.0861077517, -24.0270462386, -4.15059590987, -3.92373950824, -59.3656430833, 19.7314181435, -96.4668701748};
test_label[1455] = '{19.7314181435};
test_output[1455] = '{9.57749435361e-11};
############ END DEBUG ############*/
test_input[11648:11655] = '{32'h42b976a5, 32'h40b523b6, 32'h41200486, 32'hc2bf4778, 32'hc118fa93, 32'h409f5392, 32'hc2a40c9e, 32'hc252eb5f};
test_label[1456] = '{32'h41200486};
test_output[1456] = '{32'h42a57614};
/*############ DEBUG ############
test_input[11648:11655] = '{92.7317241731, 5.66060931736, 10.0011040107, -95.6395861969, -9.56117574866, 4.97895129165, -82.0246448813, -52.7298544851};
test_label[1456] = '{10.0011040107};
test_output[1456] = '{82.7306201624};
############ END DEBUG ############*/
test_input[11656:11663] = '{32'hbffc8c4c, 32'h419cce8b, 32'hc23f001f, 32'h416f0afe, 32'hc2a3fb85, 32'h42b76564, 32'hc24afc92, 32'hc276b051};
test_label[1457] = '{32'hbffc8c4c};
test_output[1457] = '{32'h42bb5795};
/*############ DEBUG ############
test_input[11656:11663] = '{-1.97303146142, 19.6008501766, -47.7501170788, 14.9401834927, -81.9912525179, 91.698026415, -50.7466506805, -61.6721825476};
test_label[1457] = '{-1.97303146142};
test_output[1457] = '{93.6710578764};
############ END DEBUG ############*/
test_input[11664:11671] = '{32'hc29cd4c3, 32'h41470752, 32'hc2beae83, 32'h425e9c89, 32'h404bb5c9, 32'hc294afd1, 32'h42ba2663, 32'hc1975aba};
test_label[1458] = '{32'h404bb5c9};
test_output[1458] = '{32'h42b3c8b5};
/*############ DEBUG ############
test_input[11664:11671] = '{-78.4155505826, 12.4392868597, -95.3408430175, 55.6528654616, 3.18297038348, -74.3433901815, 93.0749735987, -18.9192992397};
test_label[1458] = '{3.18297038348};
test_output[1458] = '{89.8920032152};
############ END DEBUG ############*/
test_input[11672:11679] = '{32'h4172a326, 32'h42342aae, 32'h42b7cf54, 32'h41eb5f6e, 32'hc1d30ee3, 32'h424af887, 32'h42be5760, 32'h429979e7};
test_label[1459] = '{32'h42b7cf54};
test_output[1459] = '{32'h40536755};
/*############ DEBUG ############
test_input[11672:11679] = '{15.1648314415, 45.0416808783, 91.9049350005, 29.4215961436, -26.3822681557, 50.7427010821, 95.1706578608, 76.7380942599};
test_label[1459] = '{91.9049350005};
test_output[1459] = '{3.30318177619};
############ END DEBUG ############*/
test_input[11680:11687] = '{32'hc23b795a, 32'hc29fa5d8, 32'h429d69c7, 32'hc0e764eb, 32'h42b2c414, 32'hc23fb2ee, 32'hc29aa14b, 32'hc2a2338e};
test_label[1460] = '{32'hc23fb2ee};
test_output[1460] = '{32'h43094ec7};
/*############ DEBUG ############
test_input[11680:11687] = '{-46.8685055416, -79.8239135241, 78.7065956019, -7.23106928322, 89.38296614, -47.9247374401, -77.3150283591, -81.1006922772};
test_label[1460] = '{-47.9247374401};
test_output[1460] = '{137.307726664};
############ END DEBUG ############*/
test_input[11688:11695] = '{32'hc2365521, 32'hc167fbb4, 32'h42802623, 32'hc16b9adf, 32'h413efab6, 32'h41fbd784, 32'h42631f44, 32'h41c9fed7};
test_label[1461] = '{32'h41fbd784};
test_output[1461] = '{32'h42026136};
/*############ DEBUG ############
test_input[11688:11695] = '{-45.5831336334, -14.4989513072, 64.0744865124, -14.7253099058, 11.9362085492, 31.4802326758, 56.7805328998, 25.2494336366};
test_label[1461] = '{31.4802326758};
test_output[1461] = '{32.5949332415};
############ END DEBUG ############*/
test_input[11696:11703] = '{32'h4200b073, 32'h4280117c, 32'hc2c4f10d, 32'h3ff1cffc, 32'h41bb80a3, 32'h426db0de, 32'h41dd172e, 32'hc21cef4a};
test_label[1462] = '{32'h41bb80a3};
test_output[1462] = '{32'h42226cc7};
/*############ DEBUG ############
test_input[11696:11703] = '{32.172312201, 64.0341503427, -98.470798897, 1.88915962242, 23.4378117662, 59.4227206821, 27.636318938, -39.2336807689};
test_label[1462] = '{23.4378117662};
test_output[1462] = '{40.606227124};
############ END DEBUG ############*/
test_input[11704:11711] = '{32'h42773d84, 32'h42b798b5, 32'h42c44039, 32'hc2951622, 32'hc2b99c6e, 32'hc0e86c86, 32'hc1c23fe4, 32'h42a98e3e};
test_label[1463] = '{32'hc2951622};
test_output[1463] = '{32'h432caba3};
/*############ DEBUG ############
test_input[11704:11711] = '{61.8100745971, 91.7982568397, 98.1254362965, -74.5432299211, -92.8055294611, -7.26324746615, -24.2811970994, 84.7778152782};
test_label[1463] = '{-74.5432299211};
test_output[1463] = '{172.670453284};
############ END DEBUG ############*/
test_input[11712:11719] = '{32'h42af2c3c, 32'h429b8ae3, 32'hc2a36545, 32'hc15119ec, 32'h41a1e206, 32'h42bbe4c7, 32'hc28d8c03, 32'h42863d5e};
test_label[1464] = '{32'h42863d5e};
test_output[1464] = '{32'h41d6a12a};
/*############ DEBUG ############
test_input[11712:11719] = '{87.586395581, 77.7712662764, -81.6977947225, -13.0688284092, 20.2353621825, 93.9468272883, -70.7734593964, 67.1198610221};
test_label[1464] = '{67.1198610221};
test_output[1464] = '{26.8286934884};
############ END DEBUG ############*/
test_input[11720:11727] = '{32'h4275e21e, 32'hc2b3c862, 32'h429ee330, 32'hc242946e, 32'h424014f4, 32'h42ac031d, 32'hc284752f, 32'h4294364a};
test_label[1465] = '{32'h42ac031d};
test_output[1465] = '{32'h3ab9e757};
/*############ DEBUG ############
test_input[11720:11727] = '{61.4708163085, -89.8913700227, 79.4437242819, -48.6449525848, 48.0204614388, 86.0060839599, -66.2288779247, 74.1060358992};
test_label[1465] = '{86.0060839599};
test_output[1465] = '{0.0014183324063};
############ END DEBUG ############*/
test_input[11728:11735] = '{32'hc2bb42b7, 32'h41a93049, 32'hc2bccea2, 32'hc12533b5, 32'hc2001e93, 32'hc18cee56, 32'hc2448798, 32'h4196ba4d};
test_label[1466] = '{32'hc2bccea2};
test_output[1466] = '{32'h42e74b45};
/*############ DEBUG ############
test_input[11728:11735] = '{-93.6303026767, 21.1485762968, -94.4035821178, -10.3251237515, -32.0298557377, -17.6163753419, -49.1324160919, 18.8409679381};
test_label[1466] = '{-94.4035821178};
test_output[1466] = '{115.647012975};
############ END DEBUG ############*/
test_input[11736:11743] = '{32'hc26ea08a, 32'h3f1a578e, 32'hc1e30763, 32'h42baf21e, 32'hc2c2f78b, 32'hc16eca08, 32'hc168ab92, 32'hc240a2a2};
test_label[1467] = '{32'hc2c2f78b};
test_output[1467] = '{32'h433ef4d5};
/*############ DEBUG ############
test_input[11736:11743] = '{-59.6567771956, 0.602898483266, -28.3786061709, 93.4728825905, -97.4834853803, -14.9243235882, -14.5418873428, -48.1588218261};
test_label[1467] = '{-97.4834853803};
test_output[1467] = '{190.956367971};
############ END DEBUG ############*/
test_input[11744:11751] = '{32'h4267c70e, 32'hc1042b6f, 32'hc2b46b10, 32'hc2498d25, 32'h42ade906, 32'h423ad250, 32'hc2991fb2, 32'h42354d81};
test_label[1468] = '{32'hc2b46b10};
test_output[1468] = '{32'h43312a0b};
/*############ DEBUG ############
test_input[11744:11751] = '{57.9443907778, -8.26060362771, -90.2091083282, -50.3878364831, 86.955127511, 46.705384391, -76.5619049177, 45.3256876835};
test_label[1468] = '{-90.2091083282};
test_output[1468] = '{177.164235839};
############ END DEBUG ############*/
test_input[11752:11759] = '{32'hc209d158, 32'hc294fc53, 32'hc2802415, 32'h42bd8e87, 32'h421ff844, 32'hc1255e14, 32'hc2c02aba, 32'h42bff14d};
test_label[1469] = '{32'hc2802415};
test_output[1469] = '{32'h43204e83};
/*############ DEBUG ############
test_input[11752:11759] = '{-34.4544359816, -74.4928215082, -64.0704712618, 94.778372678, 39.9924459422, -10.3354680227, -96.0834488123, 95.9712870341};
test_label[1469] = '{-64.0704712618};
test_output[1469] = '{160.306685386};
############ END DEBUG ############*/
test_input[11760:11767] = '{32'hc2b57a96, 32'hc13ead83, 32'hc2ab3f9a, 32'hbe9949a1, 32'hc1693c6d, 32'hc203975e, 32'h4271a3ad, 32'hc0bd78d5};
test_label[1470] = '{32'hc2b57a96};
test_output[1470] = '{32'h43172636};
/*############ DEBUG ############
test_input[11760:11767] = '{-90.73942439, -11.9173608042, -85.6242222341, -0.299389879147, -14.5772521235, -32.897819185, 60.4098383316, -5.92099980835};
test_label[1470] = '{-90.73942439};
test_output[1470] = '{151.149262722};
############ END DEBUG ############*/
test_input[11768:11775] = '{32'h426d67fd, 32'h42a48c94, 32'h4104f8ce, 32'hc127a3b3, 32'hc28b02f3, 32'h42bf5152, 32'h427f448f, 32'h425d6319};
test_label[1471] = '{32'hc127a3b3};
test_output[1471] = '{32'h42d445c9};
/*############ DEBUG ############
test_input[11768:11775] = '{59.3515515203, 82.2745701134, 8.31074336644, -10.4774654307, -69.5057598205, 95.6588293116, 63.8169529661, 55.3467738923};
test_label[1471] = '{-10.4774654307};
test_output[1471] = '{106.136296281};
############ END DEBUG ############*/
test_input[11776:11783] = '{32'hc2292455, 32'h42b8eb76, 32'h3fd80c20, 32'hc045faf9, 32'hc1cf6d1b, 32'h4178e065, 32'hbf8a5029, 32'h421053f6};
test_label[1472] = '{32'hc1cf6d1b};
test_output[1472] = '{32'h42ecc6bc};
/*############ DEBUG ############
test_input[11776:11783] = '{-42.2854789149, 92.4598814305, 1.68787006424, -3.09344324213, -25.9282746618, 15.5547835795, -1.08057129691, 36.0819943635};
test_label[1472] = '{-25.9282746618};
test_output[1472] = '{118.388156092};
############ END DEBUG ############*/
test_input[11784:11791] = '{32'h42c021ba, 32'hbf080e62, 32'hc1248503, 32'hc25fb029, 32'h42b3d5cf, 32'h42784fa3, 32'hc16c194c, 32'h42766199};
test_label[1473] = '{32'h42b3d5cf};
test_output[1473] = '{32'h40c4d034};
/*############ DEBUG ############
test_input[11784:11791] = '{96.0658732312, -0.53146949069, -10.2824731195, -55.9220315985, 89.9175927728, 62.0777711638, -14.7561758127, 61.5953085752};
test_label[1473] = '{89.9175927728};
test_output[1473] = '{6.15041533149};
############ END DEBUG ############*/
test_input[11792:11799] = '{32'h4201086e, 32'h4295f61b, 32'hc2b702e6, 32'hc2b339c8, 32'hc2b24656, 32'h41b058e7, 32'hc243f7e0, 32'hc1dbc05c};
test_label[1474] = '{32'hc2b339c8};
test_output[1474] = '{32'h432497f2};
/*############ DEBUG ############
test_input[11792:11799] = '{32.2582312066, 74.9806776163, -91.5056631353, -89.6128572755, -89.1373762515, 22.043410215, -48.992065132, -27.4689251699};
test_label[1474] = '{-89.6128572755};
test_output[1474] = '{164.593534892};
############ END DEBUG ############*/
test_input[11800:11807] = '{32'h404f3c7f, 32'hc1be0d5c, 32'h4220dd0d, 32'hc284bebb, 32'h424d7184, 32'hc1dd2eef, 32'h4197b445, 32'hc20c01df};
test_label[1475] = '{32'h424d7184};
test_output[1475] = '{32'h37726359};
/*############ DEBUG ############
test_input[11800:11807] = '{3.23806749904, -23.7565227241, 40.2158693018, -66.3725188108, 51.3608543372, -27.6479159246, 18.9630224924, -35.0018256833};
test_label[1475] = '{51.3608543372};
test_output[1475] = '{1.44474553602e-05};
############ END DEBUG ############*/
test_input[11808:11815] = '{32'hc292e1cf, 32'hc225cc0b, 32'h42af9cf4, 32'h418f9965, 32'hc2459026, 32'hbefa8acf, 32'h40fa9f1b, 32'hc29114fe};
test_label[1476] = '{32'hc292e1cf};
test_output[1476] = '{32'h43213f62};
/*############ DEBUG ############
test_input[11808:11815] = '{-73.4410346683, -41.449259021, 87.806550351, 17.9499003229, -49.39076884, -0.489340279315, 7.83192223249, -72.5410018326};
test_label[1476] = '{-73.4410346683};
test_output[1476] = '{161.247585019};
############ END DEBUG ############*/
test_input[11816:11823] = '{32'hc2557f15, 32'hc2189e41, 32'h423ae8eb, 32'hc2b222a7, 32'hc28bdf2d, 32'hc24b38d9, 32'hc28adf14, 32'h429eae8d};
test_label[1477] = '{32'h429eae8d};
test_output[1477] = '{32'h27f80000};
/*############ DEBUG ############
test_input[11816:11823] = '{-53.3741047052, -38.1545445285, 46.7274570556, -89.0676796057, -69.9358886758, -50.8055156833, -69.435696218, 79.3409182615};
test_label[1477] = '{79.3409182615};
test_output[1477] = '{6.88338275268e-15};
############ END DEBUG ############*/
test_input[11824:11831] = '{32'hbf6ebe70, 32'h429c5df0, 32'h428110ad, 32'hc1c76b2b, 32'h40fbea9d, 32'hc2a13da3, 32'h42999627, 32'hc2a7c3dd};
test_label[1478] = '{32'h42999627};
test_output[1478] = '{32'h3fce68a4};
/*############ DEBUG ############
test_input[11824:11831] = '{-0.932593369842, 78.1834718051, 64.5325684799, -24.9273273079, 7.87238923157, -80.6203819623, 76.7932670049, -83.8825450272};
test_label[1478] = '{76.7932670049};
test_output[1478] = '{1.61256842994};
############ END DEBUG ############*/
test_input[11832:11839] = '{32'h42bd6f76, 32'hc2b6b9cc, 32'hc182b9a5, 32'h42b3c903, 32'hc291412d, 32'hc268b2fb, 32'hc028b420, 32'hc21f8b4a};
test_label[1479] = '{32'hc291412d};
test_output[1479] = '{32'h43275a5e};
/*############ DEBUG ############
test_input[11832:11839] = '{94.7177008677, -91.3628825378, -16.340647142, 89.892598207, -72.6272982008, -58.1747849818, -2.63599403642, -39.8860261798};
test_label[1479] = '{-72.6272982008};
test_output[1479] = '{167.352992764};
############ END DEBUG ############*/
test_input[11840:11847] = '{32'hc0cb2ebe, 32'hc29fb9fc, 32'h41412197, 32'h428565fd, 32'hc1a839c8, 32'hc1fffa93, 32'h4204a06f, 32'hc242965a};
test_label[1480] = '{32'hc0cb2ebe};
test_output[1480] = '{32'h429218e9};
/*############ DEBUG ############
test_input[11840:11847] = '{-6.34945577094, -79.8632493863, 12.0707002354, 66.6991978131, -21.0282126503, -31.9973501524, 33.1566738742, -48.6468272754};
test_label[1480] = '{-6.34945577094};
test_output[1480] = '{73.048653584};
############ END DEBUG ############*/
test_input[11848:11855] = '{32'h420e72a3, 32'h42ab8864, 32'hc1b9ff9c, 32'h42845b4f, 32'h427628da, 32'hc19ffe70, 32'hc232c6a6, 32'hc2c296da};
test_label[1481] = '{32'hc1b9ff9c};
test_output[1481] = '{32'h42da084b};
/*############ DEBUG ############
test_input[11848:11855] = '{35.6119484624, 85.7663852892, -23.2498083452, 66.1783345148, 61.5398924844, -19.9992375096, -44.6939921412, -97.2946312906};
test_label[1481] = '{-23.2498083452};
test_output[1481] = '{109.016193638};
############ END DEBUG ############*/
test_input[11856:11863] = '{32'h4264999b, 32'hc2a234f3, 32'hc29e8b6c, 32'hc190ebf4, 32'hc216fffc, 32'hc13c7d79, 32'h4218ae06, 32'hc2858818};
test_label[1482] = '{32'hc190ebf4};
test_output[1482] = '{32'h429687ca};
/*############ DEBUG ############
test_input[11856:11863] = '{57.150003622, -81.1034198989, -79.2723100905, -18.1152121522, -37.7499851775, -11.7806325743, 38.1699457156, -66.7658069309};
test_label[1482] = '{-18.1152121522};
test_output[1482] = '{75.2652157799};
############ END DEBUG ############*/
test_input[11864:11871] = '{32'hc2058b44, 32'h41098c0c, 32'h42962fb5, 32'hc284c0f3, 32'hc2a3bc03, 32'h429aa799, 32'hc144a234, 32'h42735d01};
test_label[1483] = '{32'h429aa799};
test_output[1483] = '{32'h3dd05684};
/*############ DEBUG ############
test_input[11864:11871] = '{-33.3860031762, 8.59669142544, 75.0931771685, -66.3768510605, -81.8672110062, 77.3273403266, -12.2896004505, 60.8408231221};
test_label[1483] = '{77.3273403266};
test_output[1483] = '{0.101727519117};
############ END DEBUG ############*/
test_input[11872:11879] = '{32'hbe217ba7, 32'hc2686dbe, 32'hc1ad23f9, 32'h4205fdc1, 32'hc0e6a17b, 32'h428601c9, 32'h3f38cfc2, 32'h42a1f768};
test_label[1484] = '{32'h4205fdc1};
test_output[1484] = '{32'h423df10f};
/*############ DEBUG ############
test_input[11872:11879] = '{-0.157698253558, -58.1071685491, -21.6425643037, 33.4978051178, -7.20721174725, 67.0034899674, 0.721920128688, 80.9832125801};
test_label[1484] = '{33.4978051178};
test_output[1484] = '{47.4854083108};
############ END DEBUG ############*/
test_input[11880:11887] = '{32'hc07c263f, 32'h4237a060, 32'h42126102, 32'hc2183da6, 32'hc284d159, 32'h41b59e4c, 32'hc1585171, 32'hc09072f8};
test_label[1485] = '{32'hc2183da6};
test_output[1485] = '{32'h42a7ef0f};
/*############ DEBUG ############
test_input[11880:11887] = '{-3.93983426071, 45.9066149908, 36.5947334172, -38.0602027117, -66.4088830851, 22.7022934474, -13.5198828509, -4.51403447568};
test_label[1485] = '{-38.0602027117};
test_output[1485] = '{83.9669080429};
############ END DEBUG ############*/
test_input[11888:11895] = '{32'h42bcc225, 32'h428d43d2, 32'h4226d594, 32'hc1db24df, 32'h4276149c, 32'h42c43e51, 32'hc2b584cf, 32'h42783faf};
test_label[1486] = '{32'h42c43e51};
test_output[1486] = '{32'h3cbfd6d8};
/*############ DEBUG ############
test_input[11888:11895] = '{94.3791871828, 70.6324649049, 41.7085727128, -27.3930030078, 61.520124495, 98.1217110638, -90.759390798, 62.0621895823};
test_label[1486] = '{98.1217110638};
test_output[1486] = '{0.0234178747949};
############ END DEBUG ############*/
test_input[11896:11903] = '{32'h4251ae5a, 32'h420c748a, 32'h42258463, 32'h42a03ef5, 32'h412356ce, 32'hc2873d2b, 32'hc28d7277, 32'hc1bec685};
test_label[1487] = '{32'h412356ce};
test_output[1487] = '{32'h428bd41b};
/*############ DEBUG ############
test_input[11896:11903] = '{52.4202636286, 35.1138067548, 41.3792836432, 80.1229614121, 10.2086924171, -67.6194693222, -70.7235610009, -23.8469335146};
test_label[1487] = '{10.2086924171};
test_output[1487] = '{69.914268995};
############ END DEBUG ############*/
test_input[11904:11911] = '{32'hc1d63c42, 32'h42b931b9, 32'hc1c5a107, 32'hc228ca18, 32'hc28e9a35, 32'h4143a639, 32'hc27d26e0, 32'hc283f7e5};
test_label[1488] = '{32'hc1c5a107};
test_output[1488] = '{32'h42ea99fb};
/*############ DEBUG ############
test_input[11904:11911] = '{-26.7794233151, 92.5971150935, -24.7036257395, -42.1973588219, -71.301186098, 12.228081309, -63.2879627799, -65.9841703841};
test_label[1488] = '{-24.7036257395};
test_output[1488] = '{117.300740833};
############ END DEBUG ############*/
test_input[11912:11919] = '{32'h417ba81b, 32'hc0480db2, 32'hc20702db, 32'hc1acfbbd, 32'h42b48eae, 32'h42802476, 32'hc1536c57, 32'hc102acb7};
test_label[1489] = '{32'h417ba81b};
test_output[1489] = '{32'h429519ab};
/*############ DEBUG ############
test_input[11912:11919] = '{15.728541426, -3.12583589364, -33.752786726, -21.6229184968, 90.2786740107, 64.0712165473, -13.2139503605, -8.16716629937};
test_label[1489] = '{15.728541426};
test_output[1489] = '{74.5501325848};
############ END DEBUG ############*/
test_input[11920:11927] = '{32'hc161bcf3, 32'hc120a3a2, 32'hc291033a, 32'hc2b9b823, 32'h4255ac3e, 32'hc10b7d07, 32'h429178e9, 32'hc29cffa4};
test_label[1490] = '{32'hc120a3a2};
test_output[1490] = '{32'h42a58d5d};
/*############ DEBUG ############
test_input[11920:11927] = '{-14.1086304733, -10.039949327, -72.5063024588, -92.8596393856, 53.4182057433, -8.71802446454, 72.7361495348, -78.4992953553};
test_label[1490] = '{-10.039949327};
test_output[1490] = '{82.7760988659};
############ END DEBUG ############*/
test_input[11928:11935] = '{32'hc2928192, 32'hc20bc6ec, 32'hc2aa6ca9, 32'h422e75ec, 32'h41fa3f4e, 32'hc16fa603, 32'h415c3d3e, 32'h423b02d5};
test_label[1491] = '{32'h423b02d5};
test_output[1491] = '{32'h3d2df6e0};
/*############ DEBUG ############
test_input[11928:11935] = '{-73.2530674514, -34.9442607514, -85.2122239207, 43.6151571281, 31.2809113817, -14.9780297553, 13.7649521754, 46.7527661842};
test_label[1491] = '{46.7527661842};
test_output[1491] = '{0.0424717682156};
############ END DEBUG ############*/
test_input[11936:11943] = '{32'hc2a8a43a, 32'hc2828150, 32'hc18eb7de, 32'hc0d636d2, 32'h42ab0fa4, 32'hc29c2623, 32'hc2b432cd, 32'h42b0035c};
test_label[1492] = '{32'h42b0035c};
test_output[1492] = '{32'h3da5558d};
/*############ DEBUG ############
test_input[11936:11943] = '{-84.3207560136, -65.2525634023, -17.839778452, -6.69419201217, 85.5305505364, -78.0744871432, -90.0992178661, 88.0065644034};
test_label[1492] = '{88.0065644034};
test_output[1492] = '{0.0807295825686};
############ END DEBUG ############*/
test_input[11944:11951] = '{32'h427d1b3f, 32'hc25e0edc, 32'hc27a993a, 32'hc1398c0e, 32'hc28f9ee9, 32'hc28973ca, 32'h4296eba2, 32'hc28fd259};
test_label[1493] = '{32'hc28fd259};
test_output[1493] = '{32'h43135efe};
/*############ DEBUG ############
test_input[11944:11951] = '{63.2766087737, -55.5145124644, -62.649636228, -11.5966935139, -71.8103710886, -68.7261512011, 75.4602195838, -71.9108388743};
test_label[1493] = '{-71.9108388743};
test_output[1493] = '{147.371063572};
############ END DEBUG ############*/
test_input[11952:11959] = '{32'h42bee7a8, 32'h425e734a, 32'h429c0187, 32'h41fcbe89, 32'hc29a9ab1, 32'hc29c4943, 32'h4283e3c8, 32'hc2147bfa};
test_label[1494] = '{32'hc29c4943};
test_output[1494] = '{32'h432d9876};
/*############ DEBUG ############
test_input[11952:11959] = '{95.4524557687, 55.612585769, 78.0029866716, 31.5930354266, -77.3021325248, -78.1430916427, 65.9448832467, -37.1210712821};
test_label[1494] = '{-78.1430916427};
test_output[1494] = '{173.595547438};
############ END DEBUG ############*/
test_input[11960:11967] = '{32'h41007282, 32'h4264f875, 32'hc2b981a2, 32'h402408ab, 32'h4249cbd1, 32'hc28cac31, 32'h42198958, 32'hc22dbce1};
test_label[1495] = '{32'hc22dbce1};
test_output[1495] = '{32'h42c95b3e};
/*############ DEBUG ############
test_input[11960:11967] = '{8.02795590616, 57.2426345148, -92.7531881656, 2.56302904617, 50.4490382696, -70.336310999, 38.3841240824, -43.4344505576};
test_label[1495] = '{-43.4344505576};
test_output[1495] = '{100.678205381};
############ END DEBUG ############*/
test_input[11968:11975] = '{32'hc29ce3a9, 32'hc0f9accd, 32'h42b98d04, 32'h4193426b, 32'h41c48525, 32'hc0dec21d, 32'hc2b25204, 32'h42022f36};
test_label[1496] = '{32'h4193426b};
test_output[1496] = '{32'h4294bc69};
/*############ DEBUG ############
test_input[11968:11975] = '{-78.4446493659, -7.80234379732, 92.7754205227, 18.4074307388, 24.56501267, -6.9611954531, -89.1601873006, 32.5461027504};
test_label[1496] = '{18.4074307388};
test_output[1496] = '{74.367989784};
############ END DEBUG ############*/
test_input[11976:11983] = '{32'h420ed2a4, 32'h41f96714, 32'hc0a110e8, 32'h420a76bd, 32'h42c28e4b, 32'hc28d39f2, 32'h4109778d, 32'hc22c0330};
test_label[1497] = '{32'hc0a110e8};
test_output[1497] = '{32'h42cc9f5a};
/*############ DEBUG ############
test_input[11976:11983] = '{35.705704917, 31.1753302056, -5.03331365707, 34.6159567956, 97.2779190858, -70.6131736183, 8.59168720779, -43.0031110508};
test_label[1497] = '{-5.03331365707};
test_output[1497] = '{102.311232743};
############ END DEBUG ############*/
test_input[11984:11991] = '{32'h4211fd75, 32'hc1eb67ad, 32'h42c59948, 32'hc1154768, 32'h42c75c72, 32'hc2ae69f9, 32'hc1af3a7c, 32'h42a56fcf};
test_label[1498] = '{32'hc1eb67ad};
test_output[1498] = '{32'h430173ec};
/*############ DEBUG ############
test_input[11984:11991] = '{36.4975164958, -29.4256226831, 98.7993777864, -9.32993351172, 99.6805599721, -87.2069770143, -21.9035568133, 82.71837609};
test_label[1498] = '{-29.4256226831};
test_output[1498] = '{129.45281234};
############ END DEBUG ############*/
test_input[11992:11999] = '{32'h42189e4c, 32'hc0993f78, 32'h428a5f58, 32'hc22a84a6, 32'hc2822755, 32'hc22e6973, 32'hc1f2f837, 32'h421f08e2};
test_label[1499] = '{32'h421f08e2};
test_output[1499] = '{32'h41eb6b9d};
/*############ DEBUG ############
test_input[11992:11999] = '{38.1545870524, -4.78899781893, 69.1862214626, -42.6295376581, -65.0768199625, -43.6029791963, -30.3711982191, 39.7586755715};
test_label[1499] = '{39.7586755715};
test_output[1499] = '{29.4275458912};
############ END DEBUG ############*/
test_input[12000:12007] = '{32'hc156ccd4, 32'h42228ec3, 32'h41d527de, 32'h42a5fca9, 32'hc2bd92a6, 32'h41247b13, 32'hc20837cc, 32'h425142b1};
test_label[1500] = '{32'hc20837cc};
test_output[1500] = '{32'h42ea188f};
/*############ DEBUG ############
test_input[12000:12007] = '{-13.425006859, 40.6394156937, 26.6444657459, 82.9934765305, -94.7864232128, 10.2800478909, -34.0544890794, 52.3151300452};
test_label[1500] = '{-34.0544890794};
test_output[1500] = '{117.04796561};
############ END DEBUG ############*/
test_input[12008:12015] = '{32'hc144e9dc, 32'h428114d7, 32'h42630799, 32'hc156d2ff, 32'hc2368089, 32'hc28c47a1, 32'h41e9c8a2, 32'h41b1b052};
test_label[1501] = '{32'hc28c47a1};
test_output[1501] = '{32'h4306ae57};
/*############ DEBUG ############
test_input[12008:12015] = '{-12.307094172, 64.5407018715, 56.7574191601, -13.4265128568, -45.6255241133, -70.1399012014, 29.2229646655, 22.2110945443};
test_label[1501] = '{-70.1399012014};
test_output[1501] = '{134.681019628};
############ END DEBUG ############*/
test_input[12016:12023] = '{32'hc18ee711, 32'h42a34887, 32'hc296211e, 32'hc24309da, 32'h41d4d9db, 32'hc297baa9, 32'h421e7430, 32'h420dd7e6};
test_label[1502] = '{32'h421e7430};
test_output[1502] = '{32'h42281cdd};
/*############ DEBUG ############
test_input[12016:12023] = '{-17.8628246222, 81.6416528581, -75.0646789644, -48.75962215, 26.6063739972, -75.8645740415, 39.6134658655, 35.4608376333};
test_label[1502] = '{39.6134658655};
test_output[1502] = '{42.0281869927};
############ END DEBUG ############*/
test_input[12024:12031] = '{32'h41b1ed16, 32'h42ac11c8, 32'hc1986812, 32'hc2a80f8d, 32'hc2566b5f, 32'h425a42e5, 32'hc1b4d7be, 32'h418528fa};
test_label[1503] = '{32'h41b1ed16};
test_output[1503] = '{32'h427f2d05};
/*############ DEBUG ############
test_input[12024:12031] = '{22.2407645327, 86.0347306542, -19.0508152114, -84.0303747534, -53.6048538606, 54.565325393, -22.6053429479, 16.6450088774};
test_label[1503] = '{22.2407645327};
test_output[1503] = '{63.7939661215};
############ END DEBUG ############*/
test_input[12032:12039] = '{32'h41f5e9cb, 32'h41ae7b98, 32'hc0965de7, 32'h42b45ad2, 32'h425f8e03, 32'h41d3983a, 32'h400e03fa, 32'hc283c54d};
test_label[1504] = '{32'h42b45ad2};
test_output[1504] = '{32'h26b00000};
/*############ DEBUG ############
test_input[12032:12039] = '{30.73915648, 21.8103492704, -4.69896262998, 90.1773859327, 55.8886836032, 26.4493286869, 2.21899261436, -65.8853527449};
test_label[1504] = '{90.1773859327};
test_output[1504] = '{1.22124532709e-15};
############ END DEBUG ############*/
test_input[12040:12047] = '{32'hc29852f6, 32'hc1e0a925, 32'h427209ef, 32'hc2a06a00, 32'h421f9bca, 32'hc29e777a, 32'h42228ddb, 32'h42bd3b4b};
test_label[1505] = '{32'hc29852f6};
test_output[1505] = '{32'h432ac720};
/*############ DEBUG ############
test_input[12040:12047] = '{-76.162034246, -28.0825900303, 60.5097001423, -80.2070293361, 39.9021393681, -79.2333522921, 40.6385316553, 94.6158048241};
test_label[1505] = '{-76.162034246};
test_output[1505] = '{170.77783907};
############ END DEBUG ############*/
test_input[12048:12055] = '{32'h42a45c7b, 32'hc1a2e1a7, 32'h4218700b, 32'h419d23c8, 32'h3ef5b894, 32'hc245dd50, 32'hc230084a, 32'h41c4d108};
test_label[1506] = '{32'hc1a2e1a7};
test_output[1506] = '{32'h42cd14e4};
/*############ DEBUG ############
test_input[12048:12055] = '{82.1806235642, -20.3601819247, 38.1094166686, 19.6424710209, 0.479923850574, -49.4661252466, -44.0080947678, 24.6020660483};
test_label[1506] = '{-20.3601819247};
test_output[1506] = '{102.540805489};
############ END DEBUG ############*/
test_input[12056:12063] = '{32'h428db7c2, 32'hc288b1f3, 32'hc05d9b61, 32'h42bf3adc, 32'h42a3ddda, 32'h422e02d5, 32'hc12bf2d5, 32'hc20f569b};
test_label[1507] = '{32'h42bf3adc};
test_output[1507] = '{32'h35997189};
/*############ DEBUG ############
test_input[12056:12063] = '{70.8588983201, -68.3475600087, -3.4626084799, 95.6149633694, 81.9333069662, 43.5027656159, -10.746784723, -35.8345769751};
test_label[1507] = '{95.6149633694};
test_output[1507] = '{1.14324314462e-06};
############ END DEBUG ############*/
test_input[12064:12071] = '{32'h42af5557, 32'hc2684554, 32'h41fc4f94, 32'h429aed88, 32'hc2bd88d1, 32'hc1b71f51, 32'h411fce62, 32'h41146e37};
test_label[1508] = '{32'h42af5557};
test_output[1508] = '{32'h381b78ef};
/*############ DEBUG ############
test_input[12064:12071] = '{87.6666758746, -58.0677034975, 31.5388571095, 77.4639246203, -94.7672165727, -22.8902915198, 9.98788595364, 9.27690748556};
test_label[1508] = '{87.6666758746};
test_output[1508] = '{3.70675072251e-05};
############ END DEBUG ############*/
test_input[12072:12079] = '{32'h429eb088, 32'h414e5464, 32'h426d421c, 32'h4148b3eb, 32'hc20f5575, 32'hc289135f, 32'h4194d1b1, 32'hc2c129ac};
test_label[1509] = '{32'hc2c129ac};
test_output[1509] = '{32'h432fed1a};
/*############ DEBUG ############
test_input[12072:12079] = '{79.3447880012, 12.8956027331, 59.3145602318, 12.5439248433, -35.8334550227, -68.5378341111, 18.6023886381, -96.5813878228};
test_label[1509] = '{-96.5813878228};
test_output[1509] = '{175.926175826};
############ END DEBUG ############*/
test_input[12080:12087] = '{32'h41c4f8a7, 32'hc23185aa, 32'hc2514827, 32'hc0f279d0, 32'hc12d2283, 32'hc2943828, 32'hc11c3ed9, 32'hc2b3419d};
test_label[1510] = '{32'hc2514827};
test_output[1510] = '{32'h4299e23d};
/*############ DEBUG ############
test_input[12080:12087] = '{24.6214121096, -44.3805323131, -52.3204624821, -7.57736988353, -10.8209257818, -74.1096825554, -9.76534340325, -89.6281478741};
test_label[1510] = '{-52.3204624821};
test_output[1510] = '{76.9418745918};
############ END DEBUG ############*/
test_input[12088:12095] = '{32'hc24ed007, 32'h4285d7fb, 32'hc11a1f18, 32'hc277cda2, 32'h420c59cf, 32'hc275676b, 32'h428a1d17, 32'h4276a8b2};
test_label[1511] = '{32'h428a1d17};
test_output[1511] = '{32'h3de60478};
/*############ DEBUG ############
test_input[12088:12095] = '{-51.7031521724, 66.9218364859, -9.63259144026, -61.9508148606, 35.0877032582, -61.350994345, 69.0568149875, 61.6647405405};
test_label[1511] = '{69.0568149875};
test_output[1511] = '{0.112313213641};
############ END DEBUG ############*/
test_input[12096:12103] = '{32'h4291102e, 32'hc220d616, 32'h40fc1654, 32'hc08bbdc5, 32'h42b24a5d, 32'hc2a4bd84, 32'hc23a0ee2, 32'h41df0ae3};
test_label[1512] = '{32'h42b24a5d};
test_output[1512] = '{32'h3382d534};
/*############ DEBUG ############
test_input[12096:12103] = '{72.5315973667, -40.2090694548, 7.87772580156, -4.3669152361, 89.1452395222, -82.3701481429, -46.5145331475, 27.8803159467};
test_label[1512] = '{89.1452395222};
test_output[1512] = '{6.09237846523e-08};
############ END DEBUG ############*/
test_input[12104:12111] = '{32'h427ffe5f, 32'hc1f04e47, 32'hc256a407, 32'h410fa1d6, 32'h41d145f0, 32'h42b31c3b, 32'h42a51d99, 32'hc27604fc};
test_label[1513] = '{32'h41d145f0};
test_output[1513] = '{32'h427d966e};
/*############ DEBUG ############
test_input[12104:12111] = '{63.9984105767, -30.0382209695, -53.6601826648, 8.97701101709, 26.1591490239, 89.5551388686, 82.557805187, -61.5048683133};
test_label[1513] = '{26.1591490239};
test_output[1513] = '{63.3969037436};
############ END DEBUG ############*/
test_input[12112:12119] = '{32'hc22f2517, 32'h41f1ea12, 32'hc26a8ac3, 32'h42454655, 32'h42b0d6b0, 32'h42bfc417, 32'h420768b2, 32'hc1c994be};
test_label[1514] = '{32'h42bfc417};
test_output[1514] = '{32'h3a164ef4};
/*############ DEBUG ############
test_input[12112:12119] = '{-43.7862221788, 30.2392922937, -58.6355084399, 49.318682305, 88.4193151393, 95.8829883989, 33.8522408644, -25.1976283577};
test_label[1514] = '{95.8829883989};
test_output[1514] = '{0.0005733811014};
############ END DEBUG ############*/
test_input[12120:12127] = '{32'hc0d57ab3, 32'h42bfd4fc, 32'hc221432a, 32'h41fc48b9, 32'h42a95061, 32'hc299ed08, 32'hc2bf3a3b, 32'h4153d62a};
test_label[1515] = '{32'h42a95061};
test_output[1515] = '{32'h413424e8};
/*############ DEBUG ############
test_input[12120:12127] = '{-6.67122787759, 95.9159846164, -40.3155916524, 31.5355087475, 84.6569874159, -76.9629526799, -95.6137279729, 13.2397857023};
test_label[1515] = '{84.6569874159};
test_output[1515] = '{11.2590100912};
############ END DEBUG ############*/
test_input[12128:12135] = '{32'hc229b220, 32'h42a91d99, 32'h4247b21e, 32'h42a6dacf, 32'h4257388e, 32'h42a3b0dc, 32'h4204af5e, 32'hc1ce2f8a};
test_label[1516] = '{32'h42a6dacf};
test_output[1516] = '{32'h3fbac7df};
/*############ DEBUG ############
test_input[12128:12135] = '{-42.4239517955, 84.5578062899, 49.9239406778, 83.4273581984, 53.8052290348, 81.8454283826, 33.1712581346, -25.7732115671};
test_label[1516] = '{83.4273581984};
test_output[1516] = '{1.45922458943};
############ END DEBUG ############*/
test_input[12136:12143] = '{32'hc2c47277, 32'hc1738463, 32'h424b551c, 32'hbf811ddc, 32'h41b825ea, 32'h421ef9c5, 32'h422dbb07, 32'hc2997a6c};
test_label[1517] = '{32'hc1738463};
test_output[1517] = '{32'h42841b6c};
/*############ DEBUG ############
test_input[12136:12143] = '{-98.2235606984, -15.2198206931, 50.833115046, -1.00872371527, 23.0185126576, 39.743916772, 43.4326456125, -76.7391017123};
test_label[1517] = '{-15.2198206931};
test_output[1517] = '{66.0535617854};
############ END DEBUG ############*/
test_input[12144:12151] = '{32'hc2b2307c, 32'hc29af417, 32'h42ab6f4c, 32'h420c51d2, 32'h4209480b, 32'hc2946807, 32'hc2c3c363, 32'h42a5c56a};
test_label[1518] = '{32'h420c51d2};
test_output[1518] = '{32'h424ac761};
/*############ DEBUG ############
test_input[12144:12151] = '{-89.0946926637, -77.4767410665, 85.7173741806, 35.0799033887, 34.3203535846, -74.2031791987, -97.8816144782, 82.8855715743};
test_label[1518] = '{35.0799033887};
test_output[1518] = '{50.6947076323};
############ END DEBUG ############*/
test_input[12152:12159] = '{32'hc25b4faf, 32'h42926ffa, 32'h413ba631, 32'h42b0e22e, 32'h4207836b, 32'hc2763180, 32'hc2c0afe7, 32'h41a573ba};
test_label[1519] = '{32'h413ba631};
test_output[1519] = '{32'h42996d68};
/*############ DEBUG ############
test_input[12152:12159] = '{-54.8278169352, 73.2187036158, 11.7280742483, 88.4417569134, 33.8783392042, -61.548339085, -96.3435559558, 20.6815074875};
test_label[1519] = '{11.7280742483};
test_output[1519] = '{76.7136829098};
############ END DEBUG ############*/
test_input[12160:12167] = '{32'h42afade0, 32'h42bf4594, 32'h428cb292, 32'h4299852f, 32'hc1806dc2, 32'h42a32430, 32'h4296945b, 32'h4089ce37};
test_label[1520] = '{32'hc1806dc2};
test_output[1520] = '{32'h42df613b};
/*############ DEBUG ############
test_input[12160:12167] = '{87.8395993612, 95.6358976624, 70.3487705656, 76.7601252199, -16.0535927689, 81.5706809786, 75.2897556914, 4.30642258066};
test_label[1520] = '{-16.0535927689};
test_output[1520] = '{111.689902388};
############ END DEBUG ############*/
test_input[12168:12175] = '{32'h424b19a9, 32'hc23aa4cc, 32'h41754ddc, 32'hc21ae62d, 32'h421ff403, 32'h429daeac, 32'h423c3254, 32'h42789260};
test_label[1521] = '{32'hc23aa4cc};
test_output[1521] = '{32'h42fb0112};
/*############ DEBUG ############
test_input[12168:12175] = '{50.7750602672, -46.6609326404, 15.3315084646, -38.7247821715, 39.9882942017, 78.8411594306, 47.049150295, 62.1429428768};
test_label[1521] = '{-46.6609326404};
test_output[1521] = '{125.502092127};
############ END DEBUG ############*/
test_input[12176:12183] = '{32'h42a8455d, 32'h422e46f7, 32'h428cc6b9, 32'h421ec6ee, 32'hc2bda6ae, 32'h421ed685, 32'hc15871b1, 32'h41f2e685};
test_label[1522] = '{32'h42a8455d};
test_output[1522] = '{32'h358faf65};
/*############ DEBUG ############
test_input[12176:12183] = '{84.1354785357, 43.5693006899, 70.3881295708, 39.6942670984, -94.8255432628, 39.7094929333, -13.5277562939, 30.3625582158};
test_label[1522] = '{84.1354785357};
test_output[1522] = '{1.07053771296e-06};
############ END DEBUG ############*/
test_input[12184:12191] = '{32'h41dd7728, 32'h412592a6, 32'hc29acf15, 32'hc0c401e1, 32'hc23a4505, 32'hc12ac763, 32'h421ffe1c, 32'h42bcb558};
test_label[1523] = '{32'hc0c401e1};
test_output[1523] = '{32'h42c8f576};
/*############ DEBUG ############
test_input[12184:12191] = '{27.6831822231, 10.3483033168, -77.4044533833, -6.12522940314, -46.5674001948, -10.6736783319, 39.9981532665, 94.3541861292};
test_label[1523] = '{-6.12522940314};
test_output[1523] = '{100.479415532};
############ END DEBUG ############*/
test_input[12192:12199] = '{32'h42767658, 32'h421cc7fb, 32'hc21ed54e, 32'h427254ab, 32'h4201621b, 32'hc27aa511, 32'hc299814e, 32'h42acf7ca};
test_label[1524] = '{32'hc299814e};
test_output[1524] = '{32'h43233c8c};
/*############ DEBUG ############
test_input[12192:12199] = '{61.6155715142, 39.1952927459, -39.7083050656, 60.5826828937, 32.3458078023, -62.6611971094, -76.7525483235, 86.4839663274};
test_label[1524] = '{-76.7525483235};
test_output[1524] = '{163.236514651};
############ END DEBUG ############*/
test_input[12200:12207] = '{32'hc2adbb00, 32'hc2a19b72, 32'h42ba9ccf, 32'hc1d2961e, 32'h3ee93969, 32'h4258f4de, 32'hc28fe623, 32'h418b939a};
test_label[1525] = '{32'hc28fe623};
test_output[1525] = '{32'h43254179};
/*############ DEBUG ############
test_input[12200:12207] = '{-86.8652360379, -80.8036061789, 93.3062655497, -26.3232989816, 0.455516134411, 54.2391299791, -71.949485241, 17.4470712876};
test_label[1525] = '{-71.949485241};
test_output[1525] = '{165.255750791};
############ END DEBUG ############*/
test_input[12208:12215] = '{32'hc2b549f3, 32'h4297c88a, 32'hc0e1faf8, 32'hc201e487, 32'hc286115a, 32'h422fbf43, 32'h421a5fea, 32'hc20fa226};
test_label[1526] = '{32'hc2b549f3};
test_output[1526] = '{32'h4326893e};
/*############ DEBUG ############
test_input[12208:12215] = '{-90.6444288436, 75.8916798635, -7.06188586818, -32.4731702266, -67.0338928225, 43.9367784407, 38.593666252, -35.9083489737};
test_label[1526] = '{-90.6444288436};
test_output[1526] = '{166.536108707};
############ END DEBUG ############*/
test_input[12216:12223] = '{32'hc29d35b8, 32'h4208d595, 32'hc2a91926, 32'hc21643e3, 32'hc29e9c74, 32'h4200614d, 32'h42bf5fba, 32'hc18d206f};
test_label[1527] = '{32'hc29e9c74};
test_output[1527] = '{32'h432efe17};
/*############ DEBUG ############
test_input[12216:12223] = '{-78.6049172372, 34.2085778701, -84.5491155685, -37.5662962574, -79.3055731877, 32.0950194148, 95.6869621755, -17.6408363213};
test_label[1527] = '{-79.3055731877};
test_output[1527] = '{174.992535363};
############ END DEBUG ############*/
test_input[12224:12231] = '{32'h42b21820, 32'hc2419736, 32'hc2c736ff, 32'h41f11345, 32'h42b3abdd, 32'hc2b3e357, 32'h424e0c2b, 32'h40b8eb5e};
test_label[1528] = '{32'h42b3abdd};
test_output[1528] = '{32'h3ebfd3e8};
/*############ DEBUG ############
test_input[12224:12231] = '{89.0471199185, -48.3976659228, -99.6074114088, 30.1344090674, 89.8356728139, -89.9440215732, 51.5118834255, 5.778731383};
test_label[1528] = '{89.8356728139};
test_output[1528] = '{0.374663595731};
############ END DEBUG ############*/
test_input[12232:12239] = '{32'h42553b79, 32'hc125df3b, 32'h400233a7, 32'hc22f9a5e, 32'h42297fa8, 32'h429e36f7, 32'hc2b55f4f, 32'hc28a4349};
test_label[1529] = '{32'hc2b55f4f};
test_output[1529] = '{32'h4329cb23};
/*############ DEBUG ############
test_input[12232:12239] = '{53.3080789724, -10.3669992765, 2.03440266725, -43.9007509708, 42.3746644902, 79.1073552505, -90.6861499879, -69.1314147028};
test_label[1529] = '{-90.6861499879};
test_output[1529] = '{169.793505238};
############ END DEBUG ############*/
test_input[12240:12247] = '{32'h42bb74cb, 32'h4288a8cf, 32'hc16cbd89, 32'h4212bb52, 32'hc2a3712a, 32'h4274a28d, 32'hc287ca81, 32'h420d11de};
test_label[1530] = '{32'h4212bb52};
test_output[1530] = '{32'h42642e44};
/*############ DEBUG ############
test_input[12240:12247] = '{93.728111472, 68.3297051295, -14.7962734337, 36.6829299518, -81.7210237288, 61.1587408001, -67.895513592, 35.2674498281};
test_label[1530] = '{36.6829299518};
test_output[1530] = '{57.0451815202};
############ END DEBUG ############*/
test_input[12248:12255] = '{32'hc28c90fb, 32'h41ce6947, 32'h42a8ee10, 32'hc21c2aa8, 32'hc2680383, 32'h42c03953, 32'h427a3329, 32'h425720c2};
test_label[1531] = '{32'h427a3329};
test_output[1531] = '{32'h42063f80};
/*############ DEBUG ############
test_input[12248:12255] = '{-70.2831625541, 25.8014058751, 84.4649694461, -39.041656531, -58.003430711, 96.1119646612, 62.5499612908, 53.781988375};
test_label[1531] = '{62.5499612908};
test_output[1531] = '{33.5620121156};
############ END DEBUG ############*/
test_input[12256:12263] = '{32'hc25d1c2f, 32'hc2848077, 32'h4113a65d, 32'h429301ae, 32'h4228d840, 32'hc2b21314, 32'h42c67e3d, 32'hc2789386};
test_label[1532] = '{32'h42c67e3d};
test_output[1532] = '{32'h2ce85f00};
/*############ DEBUG ############
test_input[12256:12263] = '{-55.2775219191, -66.2509067616, 9.22811625032, 73.5032777366, 42.2111824882, -89.0372639377, 99.2465566637, -62.1440656042};
test_label[1532] = '{99.2465566637};
test_output[1532] = '{6.60438370661e-12};
############ END DEBUG ############*/
test_input[12264:12271] = '{32'hc246e393, 32'hc2012dad, 32'hc21ac4ba, 32'hbeceddff, 32'h42487e53, 32'h42a6f1be, 32'h42aa49a3, 32'h4255d018};
test_label[1533] = '{32'hc2012dad};
test_output[1533] = '{32'h42eb38a5};
/*############ DEBUG ############
test_input[12264:12271] = '{-49.7222398055, -32.294603913, -38.6921151081, -0.404037457437, 50.1233616107, 83.472150934, 85.1438183285, 53.4532165335};
test_label[1533] = '{-32.294603913};
test_output[1533] = '{117.610637438};
############ END DEBUG ############*/
test_input[12272:12279] = '{32'h4137178f, 32'h40b8d14c, 32'h42a89b59, 32'hc2590517, 32'h42219584, 32'hc28d9b91, 32'h428be02a, 32'hc0472596};
test_label[1534] = '{32'h40b8d14c};
test_output[1534] = '{32'h429d0e44};
/*############ DEBUG ############
test_input[12272:12279] = '{11.4432513915, 5.77554917149, 84.3034110972, -54.2549706759, 40.3960129597, -70.803841896, 69.9378197616, -3.11166909306};
test_label[1534] = '{5.77554917149};
test_output[1534] = '{78.5278625026};
############ END DEBUG ############*/
test_input[12280:12287] = '{32'hc13f5baf, 32'h3f94797b, 32'hc2744ac5, 32'hc15d949c, 32'hc21196d7, 32'h4269c771, 32'hc2620528, 32'h42c1d8b5};
test_label[1535] = '{32'hc13f5baf};
test_output[1535] = '{32'h42d9c42b};
/*############ DEBUG ############
test_input[12280:12287] = '{-11.9598834505, 1.15995732944, -61.0730172649, -13.8487815024, -36.3973055211, 58.4447675622, -56.505034675, 96.923255904};
test_label[1535] = '{-11.9598834505};
test_output[1535] = '{108.883139355};
############ END DEBUG ############*/
test_input[12288:12295] = '{32'hc2228f10, 32'hc2301845, 32'hc1637b4f, 32'h423bc36c, 32'h4144d946, 32'hc2844b43, 32'hc271bca3, 32'h420c1b80};
test_label[1536] = '{32'hc1637b4f};
test_output[1536] = '{32'h4274a242};
/*############ DEBUG ############
test_input[12288:12295] = '{-40.6397078359, -44.0237018968, -14.2176046504, 46.9408432803, 12.3030456844, -66.1469965548, -60.4342137144, 35.0268552494};
test_label[1536] = '{-14.2176046504};
test_output[1536] = '{61.1584546267};
############ END DEBUG ############*/
test_input[12296:12303] = '{32'hc2aed02a, 32'h424afeff, 32'h42b98a1e, 32'hc2909f5e, 32'hc0b24226, 32'hc2a1faab, 32'hc239f502, 32'h42b69248};
test_label[1537] = '{32'hc2a1faab};
test_output[1537] = '{32'h432df6b4};
/*############ DEBUG ############
test_input[12296:12303] = '{-87.4065724367, 50.7490213625, 92.7697605347, -72.3112663205, -5.57057482908, -80.9895891534, -46.489264765, 91.2857070184};
test_label[1537] = '{-80.9895891534};
test_output[1537] = '{173.963691039};
############ END DEBUG ############*/
test_input[12304:12311] = '{32'h422d27a5, 32'h41a8cfa4, 32'hc1875454, 32'hc1ef800f, 32'hc215015d, 32'h424b8bb6, 32'h42819f07, 32'h42c60250};
test_label[1538] = '{32'h424b8bb6};
test_output[1538] = '{32'h424078ea};
/*############ DEBUG ############
test_input[12304:12311] = '{43.2887157871, 21.1013872603, -16.916175393, -29.9375282596, -37.2513311409, 50.8864378201, 64.8105990594, 99.0045178197};
test_label[1538] = '{50.8864378201};
test_output[1538] = '{48.1180799995};
############ END DEBUG ############*/
test_input[12312:12319] = '{32'hc2c505bb, 32'h42aafcaf, 32'hc2c0253b, 32'h42bbbeba, 32'hc2bc9210, 32'hc243169f, 32'h428d1030, 32'hc2c6c45f};
test_label[1539] = '{32'hc2c6c45f};
test_output[1539] = '{32'h4341419b};
/*############ DEBUG ############
test_input[12312:12319] = '{-98.511191086, 85.4935194734, -96.0727188351, 93.8725103842, -94.2852795852, -48.7720911665, 70.5316197808, -99.3835357996};
test_label[1539] = '{-99.3835357996};
test_output[1539] = '{193.256275799};
############ END DEBUG ############*/
test_input[12320:12327] = '{32'hc166920e, 32'h42982a62, 32'hc26a754f, 32'h42686fa9, 32'hc272eeb4, 32'hc1961139, 32'hc27e121e, 32'hc2631e4c};
test_label[1540] = '{32'hc166920e};
test_output[1540] = '{32'h42b4fca4};
/*############ DEBUG ############
test_input[12320:12327] = '{-14.4106582669, 76.0827776306, -58.6145598327, 58.1090425503, -60.7331072105, -18.7584096921, -63.5176943968, -56.7795866994};
test_label[1540] = '{-14.4106582669};
test_output[1540] = '{90.4934359132};
############ END DEBUG ############*/
test_input[12328:12335] = '{32'hc27b6a23, 32'hc0cb5cd1, 32'h42a96b76, 32'hc1875eac, 32'h42c47eac, 32'h41a33f09, 32'hc26c6ac5, 32'hc298a420};
test_label[1541] = '{32'hc1875eac};
test_output[1541] = '{32'h42e65658};
/*############ DEBUG ############
test_input[12328:12335] = '{-62.8536477605, -6.35508007246, 84.7098830706, -16.9212264326, 98.2474095857, 20.4057786554, -59.1042671179, -76.3205603344};
test_label[1541] = '{-16.9212264326};
test_output[1541] = '{115.168637339};
############ END DEBUG ############*/
test_input[12336:12343] = '{32'hc1062435, 32'h42788251, 32'h428da798, 32'h42b205aa, 32'h428c6fde, 32'h42c51192, 32'h422cdd89, 32'h42520063};
test_label[1542] = '{32'h42520063};
test_output[1542] = '{32'h423822d4};
/*############ DEBUG ############
test_input[12336:12343] = '{-8.38383913083, 62.1272610092, 70.8273302271, 89.0110627897, 70.2184919222, 98.5343148908, 43.2163422347, 52.5003775355};
test_label[1542] = '{52.5003775355};
test_output[1542] = '{46.0340104841};
############ END DEBUG ############*/
test_input[12344:12351] = '{32'hc19eec2b, 32'h422c6d3b, 32'h42c0a9fe, 32'hc1b9e5ee, 32'hc29d3851, 32'h429814f4, 32'h40bcac86, 32'hc2a6b801};
test_label[1543] = '{32'h422c6d3b};
test_output[1543] = '{32'h4254e6c1};
/*############ DEBUG ############
test_input[12344:12351] = '{-19.8653159448, 43.1066687989, 96.3320151332, -23.2372708324, -78.6099964018, 76.0409237282, 5.89606008954, -83.3593805047};
test_label[1543] = '{43.1066687989};
test_output[1543] = '{53.2253463359};
############ END DEBUG ############*/
test_input[12352:12359] = '{32'hc2af547a, 32'hc2008092, 32'h42b36191, 32'hc1a64cbe, 32'h427c094b, 32'h41f8eaf6, 32'h42749afc, 32'h41a454cd};
test_label[1544] = '{32'h42749afc};
test_output[1544] = '{32'h41e4504c};
/*############ DEBUG ############
test_input[12352:12359] = '{-87.6649947863, -32.1255555309, 89.6905579006, -20.7874715434, 63.00907544, 31.1147265674, 61.1513513481, 20.5414072428};
test_label[1544] = '{61.1513513481};
test_output[1544] = '{28.5392065525};
############ END DEBUG ############*/
test_input[12360:12367] = '{32'hc0734b10, 32'hbfe053ba, 32'hc24ee909, 32'hc2c004b7, 32'h42a9957a, 32'h42100e8f, 32'h412a7109, 32'hc2b8b089};
test_label[1545] = '{32'h42a9957a};
test_output[1545] = '{32'h80000000};
/*############ DEBUG ############
test_input[12360:12367] = '{-3.80145645535, -1.75255517519, -51.7275723681, -96.0092057003, 84.7919437113, 36.0142185938, 10.6525960819, -92.3447931336};
test_label[1545] = '{84.7919437113};
test_output[1545] = '{-0.0};
############ END DEBUG ############*/
test_input[12368:12375] = '{32'hc17d0d0a, 32'h42c7e33f, 32'hc0b6b809, 32'h4277465d, 32'h427fe15d, 32'h40a3b4ab, 32'hc10f9c5f, 32'h421c950c};
test_label[1546] = '{32'h4277465d};
test_output[1546] = '{32'h42188020};
/*############ DEBUG ############
test_input[12368:12375] = '{-15.8156831418, 99.9438369002, -5.70996502854, 61.8187149463, 63.9700827932, 5.11580411471, -8.97567618678, 39.1455524101};
test_label[1546] = '{61.8187149463};
test_output[1546] = '{38.125121954};
############ END DEBUG ############*/
test_input[12376:12383] = '{32'h428e51eb, 32'hc005fb5c, 32'hc202d27b, 32'h41b08838, 32'hc21c4b36, 32'hc23ab598, 32'hc1cc15f5, 32'h410d2905};
test_label[1547] = '{32'hc202d27b};
test_output[1547] = '{32'h42cfbb29};
/*############ DEBUG ############
test_input[12376:12383] = '{71.1599977811, -2.09346666752, -32.705548077, 22.0665128222, -39.0734497831, -46.6773362705, -25.5107216579, 8.82251478716};
test_label[1547] = '{-32.705548077};
test_output[1547] = '{103.865545858};
############ END DEBUG ############*/
test_input[12384:12391] = '{32'hc2adb851, 32'h42bad46e, 32'h41219722, 32'hc2b7eabc, 32'h421f3b29, 32'h42893cc1, 32'h41ee9fd1, 32'hc2b75af6};
test_label[1548] = '{32'hc2adb851};
test_output[1548] = '{32'h43344660};
/*############ DEBUG ############
test_input[12384:12391] = '{-86.8599944122, 93.4149049283, 10.0993979922, -91.9584636352, 39.8077729034, 68.6186612968, 29.8280361672, -91.6776582367};
test_label[1548] = '{-86.8599944122};
test_output[1548] = '{180.274899341};
############ END DEBUG ############*/
test_input[12392:12399] = '{32'hc2330ec6, 32'h416a4a64, 32'hc25c976a, 32'hc29d5ba8, 32'h428db72c, 32'hc27b0745, 32'h415d57e2, 32'h415e8a87};
test_label[1549] = '{32'hc25c976a};
test_output[1549] = '{32'h42fc02e1};
/*############ DEBUG ############
test_input[12392:12399] = '{-44.7644253206, 14.6431620769, -55.1478661282, -78.6790182511, 70.8577589922, -62.7571006984, 13.8339554726, 13.908820439};
test_label[1549] = '{-55.1478661282};
test_output[1549] = '{126.00562512};
############ END DEBUG ############*/
test_input[12400:12407] = '{32'h424139a7, 32'h42a33c33, 32'h418d5cbc, 32'h4132dbe4, 32'h42b4d157, 32'hc29b4e52, 32'hc18b1c0e, 32'h4228d669};
test_label[1550] = '{32'h42b4d157};
test_output[1550] = '{32'h391f6d03};
/*############ DEBUG ############
test_input[12400:12407] = '{48.3063010078, 81.6175802459, 17.6702801309, 11.1786840736, 90.4088690657, -77.6529718037, -17.3886985709, 42.2093836823};
test_label[1550] = '{90.4088690657};
test_output[1550] = '{0.000152040315166};
############ END DEBUG ############*/
test_input[12408:12415] = '{32'h42391e9e, 32'hc2675861, 32'hc2c37304, 32'hc2ae0474, 32'hc2b8c282, 32'hc2334ed8, 32'hc257622f, 32'h425a584c};
test_label[1551] = '{32'hc2c37304};
test_output[1551] = '{32'h43184fa5};
/*############ DEBUG ############
test_input[12408:12415] = '{46.2799011402, -57.8363084124, -97.7246413915, -87.008699378, -92.3798982143, -44.8269951487, -53.8458807815, 54.5862260729};
test_label[1551] = '{-97.7246413915};
test_output[1551] = '{152.311114384};
############ END DEBUG ############*/
test_input[12416:12423] = '{32'h42a7903c, 32'hc2ba8f9a, 32'hc29e0d84, 32'h429dab54, 32'h41539edf, 32'h421c647a, 32'hc2b088fc, 32'hc2c1fa20};
test_label[1552] = '{32'hc2c1fa20};
test_output[1552] = '{32'h4334c6fe};
/*############ DEBUG ############
test_input[12416:12423] = '{83.7817114538, -93.280471988, -79.0263977581, 78.8346278716, 13.2262866466, 39.0981222707, -88.2675477018, -96.9885248488};
test_label[1552] = '{-96.9885248488};
test_output[1552] = '{180.777315285};
############ END DEBUG ############*/
test_input[12424:12431] = '{32'h42281904, 32'hc245659c, 32'h42bab801, 32'h4287fdcb, 32'h4278e101, 32'hc1f0e1e3, 32'hc226f783, 32'h42a51b68};
test_label[1553] = '{32'hc226f783};
test_output[1553] = '{32'h430719e2};
/*############ DEBUG ############
test_input[12424:12431] = '{42.0244308718, -49.3492260141, 93.3593805151, 67.9956860842, 62.2197305505, -30.1102963359, -41.7417109726, 82.5535307687};
test_label[1553] = '{-41.7417109726};
test_output[1553] = '{135.101111768};
############ END DEBUG ############*/
test_input[12432:12439] = '{32'h42639be0, 32'hc2b335db, 32'h426530fc, 32'h421b70e0, 32'h423a208a, 32'h4280b1ae, 32'h41fada51, 32'h429600f1};
test_label[1554] = '{32'h41fada51};
test_output[1554] = '{32'h422e94bf};
/*############ DEBUG ############
test_input[12432:12439] = '{56.9022208318, -89.6051860545, 57.2978374375, 38.8602284674, 46.5317770668, 64.3470340075, 31.3565988581, 75.0018360689};
test_label[1554] = '{31.3565988581};
test_output[1554] = '{43.6452608321};
############ END DEBUG ############*/
test_input[12440:12447] = '{32'h42c03d51, 32'h4201d23e, 32'hc20c8892, 32'hc138bef7, 32'h4140975f, 32'hc289c783, 32'h42713781, 32'h41ddbc15};
test_label[1555] = '{32'h41ddbc15};
test_output[1555] = '{32'h4288ce4c};
/*############ DEBUG ############
test_input[12440:12447] = '{96.1197598196, 32.4553146336, -35.1333704966, -11.5466223752, 12.0369554549, -68.8896713404, 60.3042042849, 27.7168375385};
test_label[1555] = '{27.7168375385};
test_output[1555] = '{68.4029222811};
############ END DEBUG ############*/
test_input[12448:12455] = '{32'hc282a6dd, 32'h41300ba5, 32'hc285eeda, 32'hc2803a5d, 32'h4037ec0c, 32'hc29d7d9e, 32'h41764766, 32'h423a8b1d};
test_label[1556] = '{32'h4037ec0c};
test_output[1556] = '{32'h422f0c5c};
/*############ DEBUG ############
test_input[12448:12455] = '{-65.3259066743, 11.0028427783, -66.9665066354, -64.1139874466, 2.87378214373, -78.7453498243, 15.3924315952, 46.6358536292};
test_label[1556] = '{2.87378214373};
test_output[1556] = '{43.7620714855};
############ END DEBUG ############*/
test_input[12456:12463] = '{32'hc25be092, 32'h42a47a86, 32'h40f72459, 32'hc2790102, 32'hc198fba7, 32'hc2a1aee1, 32'hc2142e7e, 32'h42889887};
test_label[1557] = '{32'hc2790102};
test_output[1557] = '{32'h43107d84};
/*############ DEBUG ############
test_input[12456:12463] = '{-54.9693062426, 82.2393028888, 7.72318706334, -62.2509847267, -19.1228765509, -80.8415609931, -37.0454017987, 68.2979020695};
test_label[1557] = '{-62.2509847267};
test_output[1557] = '{144.490288497};
############ END DEBUG ############*/
test_input[12464:12471] = '{32'hc2589e66, 32'hc2b10cec, 32'hc272ffb9, 32'h41551c70, 32'hc11110e2, 32'hc2c5c719, 32'hc27e757d, 32'hc1d36bd5};
test_label[1558] = '{32'hc27e757d};
test_output[1558] = '{32'h4299de4c};
/*############ DEBUG ############
test_input[12464:12471] = '{-54.1546859263, -88.5252389077, -60.7497307757, 13.3194424051, -9.06662180722, -98.8888654577, -63.6147328777, -26.4276528344};
test_label[1558] = '{-63.6147328777};
test_output[1558] = '{76.934175283};
############ END DEBUG ############*/
test_input[12472:12479] = '{32'hc298b011, 32'h428e7f18, 32'hc232d5d5, 32'h41498532, 32'hc27206c1, 32'hc262397a, 32'h4227eca0, 32'hc2207b1e};
test_label[1559] = '{32'h4227eca0};
test_output[1559] = '{32'h41ea2320};
/*############ DEBUG ############
test_input[12472:12479] = '{-76.3438764047, 71.2482286674, -44.7088203765, 12.5950182505, -60.5065959733, -56.5561312875, 41.9810775428, -40.1202300573};
test_label[1559] = '{41.9810775428};
test_output[1559] = '{29.2671511246};
############ END DEBUG ############*/
test_input[12480:12487] = '{32'hc261aafb, 32'h42c0f476, 32'hc23e56b0, 32'hc28eee6d, 32'hc1d7df8f, 32'h429f9abd, 32'h421149b4, 32'h4263b5f9};
test_label[1560] = '{32'hc1d7df8f};
test_output[1560] = '{32'h42f6ec5a};
/*############ DEBUG ############
test_input[12480:12487] = '{-56.4169727838, 96.4774646712, -47.5846541182, -71.4656746935, -26.9841594684, 79.8022224088, 36.3219753336, 56.9277095184};
test_label[1560] = '{-26.9841594684};
test_output[1560] = '{123.461624197};
############ END DEBUG ############*/
test_input[12488:12495] = '{32'hc208025e, 32'hc19e084b, 32'hc2c3e8c1, 32'h41978bdd, 32'h41ba683f, 32'h41734443, 32'hc28560b4, 32'hc28ad0a2};
test_label[1561] = '{32'h41734443};
test_output[1561] = '{32'h4101c199};
/*############ DEBUG ############
test_input[12488:12495] = '{-34.002310127, -19.7540487417, -97.9545960788, 18.9432931922, 23.3009022332, 15.2041650892, -66.6888726333, -69.4074830557};
test_label[1561] = '{15.2041650892};
test_output[1561] = '{8.10976541428};
############ END DEBUG ############*/
test_input[12496:12503] = '{32'h42b47428, 32'hc2b6dc65, 32'hc16ae832, 32'h42870a12, 32'hc230b48f, 32'h425fffac, 32'hc2b7776f, 32'hc1ac4aed};
test_label[1562] = '{32'hc16ae832};
test_output[1562] = '{32'h42d1d12e};
/*############ DEBUG ############
test_input[12496:12503] = '{90.226866918, -91.4304595001, -14.681688777, 67.519668919, -44.1763256085, 55.9996791403, -91.7332722439, -21.5365840488};
test_label[1562] = '{-14.681688777};
test_output[1562] = '{104.908555695};
############ END DEBUG ############*/
test_input[12504:12511] = '{32'h42398698, 32'h42c017d3, 32'hc22fd354, 32'h42af4137, 32'hc250e62d, 32'hc2ad51dc, 32'hc04f6994, 32'hc2b5ca57};
test_label[1563] = '{32'hc04f6994};
test_output[1563] = '{32'h42c6933d};
/*############ DEBUG ############
test_input[12504:12511] = '{46.3814403144, 96.0465315794, -43.9563735064, 87.6273764499, -52.2247791734, -86.6598822426, -3.24081891879, -90.8951984292};
test_label[1563] = '{-3.24081891879};
test_output[1563] = '{99.2875710748};
############ END DEBUG ############*/
test_input[12512:12519] = '{32'hc1373d91, 32'h41dab4ad, 32'h42c11c4a, 32'hc2c539b0, 32'h416e5573, 32'hc096652b, 32'hc2bb43b6, 32'hc2c780bd};
test_label[1564] = '{32'hc1373d91};
test_output[1564] = '{32'h42d803fc};
/*############ DEBUG ############
test_input[12512:12519] = '{-11.4525306376, 27.3382198327, 96.5552546726, -98.6126740968, 14.8958615554, -4.69984953496, -93.6322506097, -99.7514387594};
test_label[1564] = '{-11.4525306376};
test_output[1564] = '{108.00778531};
############ END DEBUG ############*/
test_input[12520:12527] = '{32'hc201099a, 32'h40d119b4, 32'h428feace, 32'h3f0f6c29, 32'h42bb0c54, 32'hc2262433, 32'h41ad4a51, 32'h41a9b991};
test_label[1565] = '{32'h3f0f6c29};
test_output[1565] = '{32'h42b9ed7c};
/*############ DEBUG ############
test_input[12520:12527] = '{-32.2593746475, 6.53438780663, 71.9586030014, 0.560244136969, 93.5240796645, -41.5353523389, 21.6612866548, 21.2156085109};
test_label[1565] = '{0.560244136969};
test_output[1565] = '{92.9638355279};
############ END DEBUG ############*/
test_input[12528:12535] = '{32'h42c453ea, 32'h40d65f03, 32'h41aaade8, 32'hc1febf60, 32'h4056d853, 32'h429492e4, 32'h416e2250, 32'h41f46b74};
test_label[1566] = '{32'h41aaade8};
test_output[1566] = '{32'h4299a870};
/*############ DEBUG ############
test_input[12528:12535] = '{98.1638957571, 6.69909800026, 21.3349157727, -31.8434454418, 3.35695348135, 74.2868948406, 14.8833770208, 30.5524668292};
test_label[1566] = '{21.3349157727};
test_output[1566] = '{76.8289799844};
############ END DEBUG ############*/
test_input[12536:12543] = '{32'h4294f185, 32'h421069ee, 32'hc2603482, 32'h4097439a, 32'hc28b5719, 32'hc2bbab7f, 32'hc26392ad, 32'hc17b5977};
test_label[1567] = '{32'h4294f185};
test_output[1567] = '{32'h80000000};
/*############ DEBUG ############
test_input[12536:12543] = '{74.4717205915, 36.1034462691, -56.0512756607, 4.72700220615, -69.6701149376, -93.8349503194, -56.8932374443, -15.7093418485};
test_label[1567] = '{74.4717205915};
test_output[1567] = '{-0.0};
############ END DEBUG ############*/
test_input[12544:12551] = '{32'hc25125cb, 32'h40aa9964, 32'hc289ca6a, 32'hc20a44bb, 32'h419be1fa, 32'h4200bc38, 32'h425afe10, 32'hc297f8f1};
test_label[1568] = '{32'h40aa9964};
test_output[1568] = '{32'h4245aae4};
/*############ DEBUG ############
test_input[12544:12551] = '{-52.2869066744, 5.3312245127, -68.8953415797, -34.5671211716, 19.4853396277, 32.1838064121, 54.7481081177, -75.9862144123};
test_label[1568] = '{5.3312245127};
test_output[1568] = '{49.4168836051};
############ END DEBUG ############*/
test_input[12552:12559] = '{32'h422aacf6, 32'h42abcd95, 32'h42291f4a, 32'hc2b04f90, 32'hc2b245f1, 32'h424fc0cf, 32'hc29e110e, 32'h42b085cc};
test_label[1569] = '{32'h424fc0cf};
test_output[1569] = '{32'h4211a731};
/*############ DEBUG ############
test_input[12552:12559] = '{42.6689089552, 85.9015252324, 42.2805562533, -88.1553989938, -89.1366056257, 51.9382914009, -79.0333073349, 88.2613209654};
test_label[1569] = '{51.9382914009};
test_output[1569] = '{36.4132719356};
############ END DEBUG ############*/
test_input[12560:12567] = '{32'hc103c67a, 32'hc02b0dca, 32'h42a6b347, 32'hc2bacd38, 32'h414a9a0e, 32'h41839750, 32'hc1b0c349, 32'h42a4227d};
test_label[1570] = '{32'hc103c67a};
test_output[1570] = '{32'h42b7a962};
/*############ DEBUG ############
test_input[12560:12567] = '{-8.2359558057, -2.67271664935, 83.3501524307, -93.4008197788, 12.6626107856, 16.4488831081, -22.095354364, 82.0673593443};
test_label[1570] = '{-8.2359558057};
test_output[1570] = '{91.8308268056};
############ END DEBUG ############*/
test_input[12568:12575] = '{32'hc1a1fa68, 32'h42becf5a, 32'hc2155529, 32'h42874e86, 32'h4219a21d, 32'hc2b6d7f3, 32'hc26ebbc4, 32'hc0356232};
test_label[1571] = '{32'hc0356232};
test_output[1571] = '{32'h42c47a6b};
/*############ DEBUG ############
test_input[12568:12575] = '{-20.2472679211, 95.4049821154, -37.3331627826, 67.6533675947, 38.4083149308, -91.4217738858, -59.683366706, -2.83411836881};
test_label[1571] = '{-2.83411836881};
test_output[1571] = '{98.2391004842};
############ END DEBUG ############*/
test_input[12576:12583] = '{32'h42acaed7, 32'h428e4849, 32'h42b95fd4, 32'hc291e4c0, 32'h41d3ec7b, 32'hc244191b, 32'h42a1a18e, 32'hc25a078e};
test_label[1572] = '{32'h42b95fd4};
test_output[1572] = '{32'h3ae6a724};
/*############ DEBUG ############
test_input[12576:12583] = '{86.3414845492, 71.1411814377, 92.6871671066, -72.9467751187, 26.4904692031, -49.0245164383, 80.8155329581, -54.5073783736};
test_label[1572] = '{92.6871671066};
test_output[1572] = '{0.00175974188331};
############ END DEBUG ############*/
test_input[12584:12591] = '{32'hc1d19156, 32'hc1c7f049, 32'h428abf40, 32'h42b51db1, 32'h42954723, 32'hc1127293, 32'h42707b4d, 32'hc210f5eb};
test_label[1573] = '{32'h42707b4d};
test_output[1573] = '{32'h41f3802a};
/*############ DEBUG ############
test_input[12584:12591] = '{-26.1959655726, -24.992327236, 69.3735372449, 90.5579907098, 74.6389413473, -9.15297241341, 60.1204101201, -36.2401537452};
test_label[1573] = '{60.1204101201};
test_output[1573] = '{30.4375807124};
############ END DEBUG ############*/
test_input[12592:12599] = '{32'hc206324c, 32'hc20c5016, 32'hc24104db, 32'h41c442bf, 32'hc289896a, 32'h420e45a7, 32'hc2bb9f8f, 32'h423361bd};
test_label[1574] = '{32'h420e45a7};
test_output[1574] = '{32'h411470bd};
/*############ DEBUG ############
test_input[12592:12599] = '{-33.5491175811, -35.0782106175, -48.2547406354, 24.5325902132, -68.7683869313, 35.5680181537, -93.8116380349, 44.8454489275};
test_label[1574] = '{35.5680181537};
test_output[1574] = '{9.27752428196};
############ END DEBUG ############*/
test_input[12600:12607] = '{32'hc1e88d92, 32'hc1087aff, 32'hc2ae4d54, 32'h40c181f7, 32'hc2303fbe, 32'hc1f7ef17, 32'hc2447680, 32'hc1c602b4};
test_label[1575] = '{32'hc2303fbe};
test_output[1575] = '{32'h42486ffd};
/*############ DEBUG ############
test_input[12600:12607] = '{-29.069125778, -8.53002874523, -87.1510304269, 6.04711478032, -44.0622478268, -30.9917439279, -49.1157240318, -24.7513204225};
test_label[1575] = '{-44.0622478268};
test_output[1575] = '{50.1093630741};
############ END DEBUG ############*/
test_input[12608:12615] = '{32'hc2a0a591, 32'hc2037485, 32'hc215594a, 32'h417f52ac, 32'h42ba8d68, 32'hc26daa81, 32'hc2c417a6, 32'hc2bc3f01};
test_label[1576] = '{32'h42ba8d68};
test_output[1576] = '{32'h80000000};
/*############ DEBUG ############
test_input[12608:12615] = '{-80.3233712345, -32.863787375, -37.3371974572, 15.9576831327, 93.2761861112, -59.416508521, -98.0461868195, -94.1230510798};
test_label[1576] = '{93.2761861112};
test_output[1576] = '{-0.0};
############ END DEBUG ############*/
test_input[12616:12623] = '{32'hc298b3b3, 32'hc219d2ad, 32'hc1e442c3, 32'h41e6f782, 32'h4211c400, 32'h42a677e7, 32'h42c4d6c7, 32'hc29d9fa6};
test_label[1577] = '{32'h42c4d6c7};
test_output[1577] = '{32'h34887369};
/*############ DEBUG ############
test_input[12616:12623] = '{-76.350973504, -38.4557366821, -28.5325986881, 28.8708534531, 36.4414054119, 83.2341807315, 98.4194846183, -78.8118157812};
test_label[1577] = '{98.4194846183};
test_output[1577] = '{2.54159449255e-07};
############ END DEBUG ############*/
test_input[12624:12631] = '{32'h42a8570e, 32'h40ae60b9, 32'hc286a77d, 32'h419844c4, 32'h429625f5, 32'h41c6720e, 32'h42b86bcc, 32'h4280b030};
test_label[1578] = '{32'h41c6720e};
test_output[1578] = '{32'h4286cf72};
/*############ DEBUG ############
test_input[12624:12631] = '{84.1700253828, 5.4493069156, -67.3271273009, 19.0335770025, 75.0741334681, 24.8056915102, 92.2105387412, 64.3441171048};
test_label[1578] = '{24.8056915102};
test_output[1578] = '{67.4051693587};
############ END DEBUG ############*/
test_input[12632:12639] = '{32'h419bf9d1, 32'hc2a6d05c, 32'h40c26fad, 32'h42361739, 32'h4221368b, 32'h4197133b, 32'h4284988f, 32'hc2bd5c9f};
test_label[1579] = '{32'h4221368b};
test_output[1579] = '{32'h41cff527};
/*############ DEBUG ############
test_input[12632:12639] = '{19.496980771, -83.4069554264, 6.07613248078, 45.5226799079, 40.303263968, 18.8843901394, 66.2979669114, -94.68089715};
test_label[1579] = '{40.303263968};
test_output[1579] = '{25.9947029444};
############ END DEBUG ############*/
test_input[12640:12647] = '{32'hc25520ca, 32'hc229a734, 32'hc2a96bba, 32'hc2c3bdb0, 32'h3f3a2abb, 32'hc2874a29, 32'h428431c4, 32'h42877787};
test_label[1580] = '{32'h42877787};
test_output[1580] = '{32'h3e362c1d};
/*############ DEBUG ############
test_input[12640:12647] = '{-53.2820196574, -42.4132859464, -84.7104067085, -97.8704833135, 0.727214521063, -67.6448457455, 66.0971990541, 67.733448162};
test_label[1580] = '{67.733448162};
test_output[1580] = '{0.177902646761};
############ END DEBUG ############*/
test_input[12648:12655] = '{32'h428fa9b7, 32'h42aed565, 32'h420a2335, 32'hc160a29a, 32'hc2be23d8, 32'hc248b775, 32'hc2b824fc, 32'h42ac174f};
test_label[1581] = '{32'hc248b775};
test_output[1581] = '{32'h4309d276};
/*############ DEBUG ############
test_input[12648:12655] = '{71.831477868, 87.4167894826, 34.5343834024, -14.0396972991, -95.0700052341, -50.1791560068, -92.0722372432, 86.0455282235};
test_label[1581] = '{-50.1791560068};
test_output[1581] = '{137.822113931};
############ END DEBUG ############*/
test_input[12656:12663] = '{32'h4087cbc3, 32'hc22545bb, 32'hc28f5423, 32'h4219403e, 32'h409eef5c, 32'h4272aa40, 32'hc2203808, 32'h421eefd8};
test_label[1582] = '{32'h4087cbc3};
test_output[1582] = '{32'h4261b0c7};
/*############ DEBUG ############
test_input[12656:12663] = '{4.24362319887, -41.3180958599, -71.6643274137, 38.3127367778, 4.96671847302, 60.6662581949, -40.0547182016, 39.7342212195};
test_label[1582] = '{4.24362319887};
test_output[1582] = '{56.4226349971};
############ END DEBUG ############*/
test_input[12664:12671] = '{32'h42907688, 32'h41f46b5b, 32'hc2acd906, 32'h42230843, 32'h415e15e8, 32'h420019a9, 32'hc2967c61, 32'hbf9b335e};
test_label[1583] = '{32'h41f46b5b};
test_output[1583] = '{32'h4226b762};
/*############ DEBUG ############
test_input[12664:12671] = '{72.2315065731, 30.5524203633, -86.4238733834, 40.7580698624, 13.8803478214, 32.0250584483, -75.2429283566, -1.21250511024};
test_label[1583] = '{30.5524203633};
test_output[1583] = '{41.6790862098};
############ END DEBUG ############*/
test_input[12672:12679] = '{32'h425d523b, 32'hc2a043b3, 32'h41393f60, 32'h41dcb2bf, 32'h41e238b8, 32'hc2284997, 32'h41be9764, 32'hc22d8b50};
test_label[1584] = '{32'hc22d8b50};
test_output[1584] = '{32'h42c56ec6};
/*############ DEBUG ############
test_input[12672:12679] = '{55.33030455, -80.132224437, 11.5779720691, 27.587279083, 28.2776951839, -42.0718661434, 23.8239203152, -43.386048977};
test_label[1584] = '{-43.386048977};
test_output[1584] = '{98.716353527};
############ END DEBUG ############*/
test_input[12680:12687] = '{32'hbfd52e56, 32'h4246cda4, 32'h41c4899b, 32'h41ea55fc, 32'h41a60491, 32'hc2377636, 32'h429c6811, 32'h413ff184};
test_label[1585] = '{32'h413ff184};
test_output[1585] = '{32'h428469e1};
/*############ DEBUG ############
test_input[12680:12687] = '{-1.66547655619, 49.7008217885, 24.5671903169, 29.2919848737, 20.7522290464, -45.8654418357, 78.2032571067, 11.9964634041};
test_label[1585] = '{11.9964634041};
test_output[1585] = '{66.2067937027};
############ END DEBUG ############*/
test_input[12688:12695] = '{32'hc23efb48, 32'h427e78ad, 32'h410f08ce, 32'hc29ac19b, 32'h423afaa7, 32'hc2800f69, 32'h4288ec0e, 32'h42c224f9};
test_label[1586] = '{32'hc2800f69};
test_output[1586] = '{32'h43211a31};
/*############ DEBUG ############
test_input[12688:12695] = '{-47.7453902297, 63.6178486658, 8.93964977392, -77.3781385716, 46.7447760712, -64.0300954657, 68.461043394, 97.072211227};
test_label[1586] = '{-64.0300954657};
test_output[1586] = '{161.102306693};
############ END DEBUG ############*/
test_input[12696:12703] = '{32'hc1b33862, 32'h42a56563, 32'h4223a64d, 32'hc28781c1, 32'h42b87a2c, 32'hc2c680a0, 32'h4148a17c, 32'h4258f8cc};
test_label[1587] = '{32'h42b87a2c};
test_output[1587] = '{32'h3896b9a3};
/*############ DEBUG ############
test_input[12696:12703] = '{-22.4025315821, 82.6980222435, 40.912404443, -67.7534291621, 92.2386191468, -99.2512196169, 12.5394246224, 54.2429661396};
test_label[1587] = '{92.2386191468};
test_output[1587] = '{7.18713502502e-05};
############ END DEBUG ############*/
test_input[12704:12711] = '{32'h42083436, 32'hc2a03f6b, 32'h4292add1, 32'h40dca5e0, 32'h428b0ba6, 32'hc22d7401, 32'h41ac5463, 32'hc096d292};
test_label[1588] = '{32'hc22d7401};
test_output[1588] = '{32'h42e972f6};
/*############ DEBUG ############
test_input[12704:12711] = '{34.050986919, -80.1238648655, 73.339485381, 6.89524851124, 69.5227484997, -43.3632861305, 21.5412039217, -4.71320437247};
test_label[1588] = '{-43.3632861305};
test_output[1588] = '{116.724532485};
############ END DEBUG ############*/
test_input[12712:12719] = '{32'hbe8543bb, 32'hc2128087, 32'hc25a681c, 32'hc282d9f6, 32'hc200f045, 32'hc29ba9f6, 32'h412bb563, 32'h4291c2b8};
test_label[1589] = '{32'hc25a681c};
test_output[1589] = '{32'h42fef6c6};
/*############ DEBUG ############
test_input[12712:12719] = '{-0.260282365219, -36.6255148639, -54.6016705888, -65.4257083256, -32.2346397847, -77.8319520685, 10.7317835019, 72.8803089299};
test_label[1589] = '{-54.6016705888};
test_output[1589] = '{127.481979519};
############ END DEBUG ############*/
test_input[12720:12727] = '{32'h428d24d0, 32'h428c15f2, 32'hc20fed3f, 32'hc0331dce, 32'h422d7da8, 32'hc29d5a68, 32'hc25952bd, 32'h42b27b68};
test_label[1590] = '{32'hc20fed3f};
test_output[1590] = '{32'h42fa7207};
/*############ DEBUG ############
test_input[12720:12727] = '{70.571901722, 70.0428599181, -35.9816845057, -2.79869414817, 43.372711909, -78.6765770224, -54.330800557, 89.2410255098};
test_label[1590] = '{-35.9816845057};
test_output[1590] = '{125.222710028};
############ END DEBUG ############*/
test_input[12728:12735] = '{32'hc22b395e, 32'h41815a9e, 32'hc1c49cb8, 32'hc2a5d46f, 32'h42be6abe, 32'hc1a57e6c, 32'h42a43190, 32'hc18861eb};
test_label[1591] = '{32'hc18861eb};
test_output[1591] = '{32'h42e08339};
/*############ DEBUG ############
test_input[12728:12735] = '{-42.8060216391, 16.1692461888, -24.5765223793, -82.9149069619, 95.2084796269, -20.6867297957, 82.0968022261, -17.0478122589};
test_label[1591] = '{-17.0478122589};
test_output[1591] = '{112.256293907};
############ END DEBUG ############*/
test_input[12736:12743] = '{32'h40ed5d9b, 32'hc29f508f, 32'h421b8687, 32'hc2842d9e, 32'hc21e3a02, 32'h42785d43, 32'hc2826296, 32'h42a496c3};
test_label[1592] = '{32'h42785d43};
test_output[1592] = '{32'h41a1a086};
/*############ DEBUG ############
test_input[12736:12743] = '{7.41767662556, -79.6573440784, 38.8813725406, -66.0890937792, -39.5566469016, 62.0910747295, -65.1925514387, 82.2944549778};
test_label[1592] = '{62.0910747295};
test_output[1592] = '{20.20338025};
############ END DEBUG ############*/
test_input[12744:12751] = '{32'hc26827dd, 32'hc28b5ebe, 32'h4279c813, 32'hc2a233e3, 32'hc2aa357d, 32'h40a33dae, 32'hc2702222, 32'h42741fe1};
test_label[1593] = '{32'hc2aa357d};
test_output[1593] = '{32'h4313c479};
/*############ DEBUG ############
test_input[12744:12751] = '{-58.038927544, -69.685040236, 62.445386546, -81.1013375515, -85.1044684389, 5.10127925845, -60.0333317625, 61.0311310598};
test_label[1593] = '{-85.1044684389};
test_output[1593] = '{147.767468508};
############ END DEBUG ############*/
test_input[12752:12759] = '{32'hc1f6cc2c, 32'hc20a9d94, 32'h42bb706f, 32'h41d1909a, 32'h41d01f29, 32'hc1acb73f, 32'h40cab488, 32'h41ded808};
test_label[1594] = '{32'h41ded808};
test_output[1594] = '{32'h4283ba6d};
/*############ DEBUG ############
test_input[12752:12759] = '{-30.8496941314, -34.6538841691, 93.7196004455, 26.1956057615, 26.0152157466, -21.589475648, 6.33453759888, 27.8554839288};
test_label[1594] = '{27.8554839288};
test_output[1594] = '{65.8641165167};
############ END DEBUG ############*/
test_input[12760:12767] = '{32'h42456498, 32'hc199fa1f, 32'hc0dd89c0, 32'hc2bc1181, 32'hc1c5ceeb, 32'h4206578e, 32'hc2083f2e, 32'h429f2827};
test_label[1595] = '{32'h4206578e};
test_output[1595] = '{32'h4237f8c0};
/*############ DEBUG ############
test_input[12760:12767] = '{49.3482346822, -19.2471302047, -6.92306538366, -94.0341896894, -24.7260349598, 33.5855030196, -34.061699721, 79.5784216304};
test_label[1595] = '{33.5855030196};
test_output[1595] = '{45.9929186108};
############ END DEBUG ############*/
test_input[12768:12775] = '{32'hc210f844, 32'hc2526e0d, 32'h417ee4f1, 32'h42b3a18a, 32'h429d2ab4, 32'h42a943c8, 32'hc2a6672a, 32'h4246e75e};
test_label[1596] = '{32'h42a943c8};
test_output[1596] = '{32'h40a60a05};
/*############ DEBUG ############
test_input[12768:12775] = '{-36.2424478366, -52.6074724331, 15.9308937005, 89.8155026952, 78.5834038768, 84.6323876276, -83.2014949517, 49.7259432136};
test_label[1596] = '{84.6323876276};
test_output[1596] = '{5.18872305769};
############ END DEBUG ############*/
test_input[12776:12783] = '{32'hc2c4227a, 32'h41e36693, 32'hc2a19cd7, 32'hc1b77887, 32'h41625a75, 32'hc2695461, 32'hc02e57ac, 32'hc25336bd};
test_label[1597] = '{32'hc02e57ac};
test_output[1597] = '{32'h41f93188};
/*############ DEBUG ############
test_input[12776:12783] = '{-98.0673337879, 28.4250841769, -80.8063292406, -22.9338514119, 14.1470838812, -58.3324003172, -2.72410107618, -52.8034556654};
test_label[1597] = '{-2.72410107618};
test_output[1597] = '{31.1491858828};
############ END DEBUG ############*/
test_input[12784:12791] = '{32'hc209cc42, 32'h427baa41, 32'hc2a8f92b, 32'hc1e0ab4e, 32'hc1df2012, 32'h41f4e190, 32'hc254038f, 32'hc25f0ee8};
test_label[1598] = '{32'hc2a8f92b};
test_output[1598] = '{32'h43136726};
/*############ DEBUG ############
test_input[12784:12791] = '{-34.4494718392, 62.9162627275, -84.4866582845, -28.083644604, -27.8906589907, 30.610137174, -53.0034738231, -55.7645586837};
test_label[1598] = '{-84.4866582845};
test_output[1598] = '{147.402921012};
############ END DEBUG ############*/
test_input[12792:12799] = '{32'h41a7d5db, 32'h422115be, 32'h42afb0de, 32'h4173b5e7, 32'hc230184e, 32'h42948f15, 32'hc2ba5bcb, 32'hc203df8b};
test_label[1599] = '{32'h422115be};
test_output[1599] = '{32'h423e4bff};
/*############ DEBUG ############
test_input[12792:12799] = '{20.9794224374, 40.2712344522, 87.8454467354, 15.2319092751, -44.0237351616, 74.2794569929, -93.1792846773, -32.9683049742};
test_label[1599] = '{40.2712344522};
test_output[1599] = '{47.5742135665};
############ END DEBUG ############*/
test_input[12800:12807] = '{32'hc2638d9e, 32'h4155b3fe, 32'h428cb072, 32'hc1f9f37a, 32'hc2ae3fb7, 32'hc11784b6, 32'hc2370a88, 32'hc20a9dcb};
test_label[1600] = '{32'hc2370a88};
test_output[1600] = '{32'h42e835b6};
/*############ DEBUG ############
test_input[12800:12807] = '{-56.8882994707, 13.3564437336, 70.3446192778, -31.243885699, -87.1244403418, -9.46989999857, -45.7602862888, -34.6540959449};
test_label[1600] = '{-45.7602862888};
test_output[1600] = '{116.104905567};
############ END DEBUG ############*/
test_input[12808:12815] = '{32'h42b28872, 32'h419d0fae, 32'hc1abaca9, 32'h41af2ab8, 32'hc273c1b5, 32'h4246b103, 32'h41b6e54e, 32'hc13b64d0};
test_label[1601] = '{32'hc13b64d0};
test_output[1601] = '{32'h42c9f50c};
/*############ DEBUG ############
test_input[12808:12815] = '{89.2664944011, 19.6326557832, -21.4593071908, 21.8958582868, -60.9391652999, 49.6728615887, 22.8619659062, -11.7121126065};
test_label[1601] = '{-11.7121126065};
test_output[1601] = '{100.978607008};
############ END DEBUG ############*/
test_input[12816:12823] = '{32'h4215deb5, 32'h428a2dac, 32'h3fbb2826, 32'h40e0946e, 32'h427ae8ac, 32'hc2b7d286, 32'hc1f272a9, 32'h42bc86fe};
test_label[1602] = '{32'h42bc86fe};
test_output[1602] = '{32'h2d4d9000};
/*############ DEBUG ############
test_input[12816:12823] = '{37.4674878675, 69.0891992254, 1.46216276791, 7.01811905104, 62.7272202578, -91.9111819718, -30.3059857651, 94.2636528438};
test_label[1602] = '{94.2636528438};
test_output[1602] = '{1.16848752896e-11};
############ END DEBUG ############*/
test_input[12824:12831] = '{32'hc2b976ce, 32'h412732ca, 32'hc1e10e47, 32'h429df9aa, 32'h42b33834, 32'hc2afdefd, 32'h426c7e01, 32'h4082511c};
test_label[1603] = '{32'hc1e10e47};
test_output[1603] = '{32'h42eb7bc9};
/*############ DEBUG ############
test_input[12824:12831] = '{-92.7320384697, 10.44989924, -28.1319709412, 78.9876234966, 89.6097733533, -87.9355218424, 59.1230504267, 4.07240086756};
test_label[1603] = '{-28.1319709412};
test_output[1603] = '{117.741768664};
############ END DEBUG ############*/
test_input[12832:12839] = '{32'hc23fc399, 32'h42c3f057, 32'h4288b359, 32'hc26a36f0, 32'hc28afaed, 32'hc29968ae, 32'h41b6bbd0, 32'hc2a0b0ad};
test_label[1604] = '{32'h42c3f057};
test_output[1604] = '{32'h2a1a4000};
/*############ DEBUG ############
test_input[12832:12839] = '{-47.9410151937, 97.9694159327, 68.3502919694, -58.5536513966, -69.4900926359, -76.7044506039, 22.8417044182, -80.3450681815};
test_label[1604] = '{97.9694159327};
test_output[1604] = '{1.37001521239e-13};
############ END DEBUG ############*/
test_input[12840:12847] = '{32'hc220db83, 32'h42b09973, 32'h4233e721, 32'hc24501bf, 32'hc2c21104, 32'hc251b494, 32'h41b32ef4, 32'hc16a06af};
test_label[1605] = '{32'h41b32ef4};
test_output[1605] = '{32'h4283cdb6};
/*############ DEBUG ############
test_input[12840:12847] = '{-40.2143685054, 88.2997059331, 44.9757128169, -49.2517061064, -97.0332329198, -52.4263475829, 22.3979255309, -14.6266320616};
test_label[1605] = '{22.3979255309};
test_output[1605] = '{65.9017804022};
############ END DEBUG ############*/
test_input[12848:12855] = '{32'hc218d69a, 32'hc20bf234, 32'h4227cd25, 32'h41c372aa, 32'h41f54ec2, 32'hc25c2165, 32'h42a5de38, 32'hc1a9f986};
test_label[1606] = '{32'hc1a9f986};
test_output[1606] = '{32'h42d05c9a};
/*############ DEBUG ############
test_input[12848:12855] = '{-38.209571468, -34.9865262795, 41.9503377593, 24.4309883369, 30.6634551076, -55.0326101859, 82.9340205236, -21.2468384392};
test_label[1606] = '{-21.2468384392};
test_output[1606] = '{104.180858963};
############ END DEBUG ############*/
test_input[12856:12863] = '{32'hc27d758c, 32'hc23b2786, 32'hc23d20c7, 32'hc2b0e04c, 32'hc2aaa8f9, 32'h41bbc938, 32'hc26ac30c, 32'h4062aebb};
test_label[1607] = '{32'hc27d758c};
test_output[1607] = '{32'h42adad14};
/*############ DEBUG ############
test_input[12856:12863] = '{-63.3647932275, -46.7885970693, -47.2820085417, -88.4380806878, -85.3300255042, 23.473250733, -58.6904749735, 3.54191465509};
test_label[1607] = '{-63.3647932275};
test_output[1607] = '{86.8380439626};
############ END DEBUG ############*/
test_input[12864:12871] = '{32'hc2441083, 32'hc21c80c9, 32'h42b4283c, 32'hc2ad973d, 32'h41f0c46d, 32'h428a0db7, 32'h41b4e417, 32'hc299e615};
test_label[1608] = '{32'h42b4283c};
test_output[1608] = '{32'h3045e814};
/*############ DEBUG ############
test_input[12864:12871] = '{-49.0161255827, -39.1257661619, 90.078586186, -86.7953855833, 30.0959101615, 69.0267883829, 22.6113724003, -76.9493818337};
test_label[1608] = '{90.078586186};
test_output[1608] = '{7.19979853773e-10};
############ END DEBUG ############*/
test_input[12872:12879] = '{32'hc257242f, 32'h4281ce6f, 32'hc21abfc7, 32'h4255da0a, 32'hc25b15d3, 32'hc2b4a72e, 32'h414717df, 32'hc20a2835};
test_label[1609] = '{32'hc25b15d3};
test_output[1609] = '{32'h42ef595a};
/*############ DEBUG ############
test_input[12872:12879] = '{-53.7853346704, 64.9031914608, -38.6872819835, 53.4629277202, -54.7713123763, -90.3265254352, 12.4433274419, -34.5392644158};
test_label[1609] = '{-54.7713123763};
test_output[1609] = '{119.674514591};
############ END DEBUG ############*/
test_input[12880:12887] = '{32'h42163c8b, 32'h4255c0f4, 32'h42973e3b, 32'hc23ef20e, 32'h42991c17, 32'hc2a9d023, 32'hc1a97795, 32'h408e789f};
test_label[1610] = '{32'hc23ef20e};
test_output[1610] = '{32'h42f93eea};
/*############ DEBUG ############
test_input[12880:12887] = '{37.5591230499, 53.4384325241, 75.6215429977, -47.7363799998, 76.5548665146, -84.9065156219, -21.1833888601, 4.45222442247};
test_label[1610] = '{-47.7363799998};
test_output[1610] = '{124.622881772};
############ END DEBUG ############*/
test_input[12888:12895] = '{32'hc2aee78d, 32'h41c010d1, 32'hc28b4c9f, 32'h42c67423, 32'hc1e945d7, 32'h42c2b1b4, 32'h423cd482, 32'h4137fb1c};
test_label[1611] = '{32'h423cd482};
test_output[1611] = '{32'h4250a539};
/*############ DEBUG ############
test_input[12888:12895] = '{-87.4522483139, 24.0082103321, -69.649651003, 99.2268318795, -29.1591020341, 97.3470767807, 47.2075257252, 11.4988061327};
test_label[1611] = '{47.2075257252};
test_output[1611] = '{52.1613502557};
############ END DEBUG ############*/
test_input[12896:12903] = '{32'h42bef0db, 32'hc1dc046d, 32'h42aea9be, 32'h42a7e2d7, 32'hc27f4b64, 32'hc155c7b9, 32'h41e80bc8, 32'hc2a669a7};
test_label[1612] = '{32'h42a7e2d7};
test_output[1612] = '{32'h4138715f};
/*############ DEBUG ############
test_input[12896:12903] = '{95.4704218291, -27.5021606508, 87.3315244171, 83.943045085, -63.8236225658, -13.3612603035, 29.005752982, -83.206354347};
test_label[1612] = '{83.943045085};
test_output[1612] = '{11.527678514};
############ END DEBUG ############*/
test_input[12904:12911] = '{32'hc295783b, 32'hc272ac88, 32'hc25f47c9, 32'hc1dfb074, 32'h424741ad, 32'hc204adbe, 32'h421a7e18, 32'hc2803945};
test_label[1613] = '{32'hc204adbe};
test_output[1613] = '{32'h42a5f7b7};
/*############ DEBUG ############
test_input[12904:12911] = '{-74.7348287047, -60.6684885808, -55.8201016602, -27.961158076, 49.8141378099, -33.1696687461, 38.623139934, -64.1118579565};
test_label[1613] = '{-33.1696687461};
test_output[1613] = '{82.9838203537};
############ END DEBUG ############*/
test_input[12912:12919] = '{32'h41fe039b, 32'hc13199d7, 32'hc28ad278, 32'h42960bf5, 32'h428a709a, 32'h423f7a05, 32'h40a1976d, 32'h42b08e70};
test_label[1614] = '{32'hc28ad278};
test_output[1614] = '{32'h431db074};
/*############ DEBUG ############
test_input[12912:12919] = '{31.7517595626, -11.1000588636, -69.4110716085, 75.0233537432, 69.2199272566, 47.8691583502, 5.04973454593, 88.2781957021};
test_label[1614] = '{-69.4110716085};
test_output[1614] = '{157.689269068};
############ END DEBUG ############*/
test_input[12920:12927] = '{32'hc2149101, 32'h4185be80, 32'hc2c21909, 32'hc238cd54, 32'hc283fc0a, 32'h4114cdcd, 32'h4297134e, 32'h407acb99};
test_label[1615] = '{32'hc238cd54};
test_output[1615] = '{32'h42f379f8};
/*############ DEBUG ############
test_input[12920:12927] = '{-37.141606407, 16.7180182795, -97.0489005587, -46.2005147022, -65.9922646895, 9.30024423472, 75.5377042615, 3.91867670678};
test_label[1615] = '{-46.2005147022};
test_output[1615] = '{121.738218964};
############ END DEBUG ############*/
test_input[12928:12935] = '{32'h42334cd0, 32'hc2a384a1, 32'hc0b87220, 32'hc2676db5, 32'hc29eb42d, 32'hc1bc0ad4, 32'hc29a56b0, 32'h429bc143};
test_label[1616] = '{32'hc29eb42d};
test_output[1616] = '{32'h431d3ab8};
/*############ DEBUG ############
test_input[12928:12935] = '{44.8250134041, -81.7590423011, -5.76393133335, -57.8571360027, -79.3519069324, -23.5052876764, -77.169314724, 77.8774659678};
test_label[1616] = '{-79.3519069324};
test_output[1616] = '{157.2293729};
############ END DEBUG ############*/
test_input[12936:12943] = '{32'h41ac0044, 32'h420371d8, 32'hc2a5ffd5, 32'h42ad6d73, 32'hc2993ac2, 32'h4264bde1, 32'hc29e5699, 32'h423ed507};
test_label[1617] = '{32'hc2a5ffd5};
test_output[1617] = '{32'h4329b6a4};
/*############ DEBUG ############
test_input[12936:12943] = '{21.5001287642, 32.8611757231, -82.9996729398, 86.7137655344, -76.6147638025, 57.1854281969, -79.1691356464, 47.7080334637};
test_label[1617] = '{-82.9996729398};
test_output[1617] = '{169.713438474};
############ END DEBUG ############*/
test_input[12944:12951] = '{32'h42b4b491, 32'h41cedd11, 32'h4071346f, 32'hc2a5d15e, 32'hc1aa8f18, 32'hc2b2ba6d, 32'hc22bb2de, 32'hc28c69bd};
test_label[1618] = '{32'h4071346f};
test_output[1618] = '{32'h42ad2aee};
/*############ DEBUG ############
test_input[12944:12951] = '{90.3526723575, 25.8579432182, 3.76882535312, -82.908919465, -21.3198707674, -89.3641100762, -42.9246731877, -70.2065173663};
test_label[1618] = '{3.76882535312};
test_output[1618] = '{86.5838470044};
############ END DEBUG ############*/
test_input[12952:12959] = '{32'h4208d8c7, 32'hbeff00c6, 32'h42b064b8, 32'hc1380eac, 32'hc04d03f9, 32'hc124ffb0, 32'hc19baaaf, 32'hc260cd80};
test_label[1619] = '{32'hbeff00c6};
test_output[1619] = '{32'h42b163b9};
/*############ DEBUG ############
test_input[12952:12959] = '{34.2116955332, -0.498052768602, 88.1967167053, -11.5035821961, -3.20336743471, -10.3124239977, -19.4583413819, -56.2006846126};
test_label[1619] = '{-0.498052768602};
test_output[1619] = '{88.6947694739};
############ END DEBUG ############*/
test_input[12960:12967] = '{32'hc1f98a3a, 32'hc2c56629, 32'hc286a37e, 32'h42208deb, 32'hc1bca4a3, 32'h42a0a52a, 32'hc2823ebe, 32'hc2430f21};
test_label[1620] = '{32'h42a0a52a};
test_output[1620] = '{32'h80000000};
/*############ DEBUG ############
test_input[12960:12967] = '{-31.1924939333, -98.6995339214, -67.3193235193, 40.1385933024, -23.5803885658, 80.3225859667, -65.1225444852, -48.7647724545};
test_label[1620] = '{80.3225859667};
test_output[1620] = '{-0.0};
############ END DEBUG ############*/
test_input[12968:12975] = '{32'h40a661fe, 32'hc28a34cb, 32'hc1e6a1de, 32'hc26ccb86, 32'hc292b173, 32'hc2c24f28, 32'hc2c6f9c1, 32'h42979586};
test_label[1621] = '{32'hc28a34cb};
test_output[1621] = '{32'h4310e528};
/*############ DEBUG ############
test_input[12968:12975] = '{5.19946187228, -69.1031099413, -28.8290364127, -59.1987522232, -73.3465811262, -97.1546057665, -99.4878021432, 75.7920379075};
test_label[1621] = '{-69.1031099413};
test_output[1621] = '{144.895147849};
############ END DEBUG ############*/
test_input[12976:12983] = '{32'h4123d256, 32'h42ad5ae3, 32'hc2b500eb, 32'h4239c16f, 32'h424fde10, 32'hc2be8575, 32'h42926c75, 32'hc2ba3cf1};
test_label[1622] = '{32'hc2b500eb};
test_output[1622] = '{32'h43312de7};
/*############ DEBUG ############
test_input[12976:12983] = '{10.2388517217, 86.6775152245, -90.5017960632, 46.4389011226, 51.9668571989, -95.2606561707, 73.2118266067, -93.1190250532};
test_label[1622] = '{-90.5017960632};
test_output[1622] = '{177.179312706};
############ END DEBUG ############*/
test_input[12984:12991] = '{32'hc24b9412, 32'hc249a1e4, 32'hc20c0808, 32'hc286a6fb, 32'h4200d7bb, 32'h4204691e, 32'h42a0cb6d, 32'h4210ee9b};
test_label[1623] = '{32'hc286a6fb};
test_output[1623] = '{32'h4313b934};
/*############ DEBUG ############
test_input[12984:12991] = '{-50.8946017894, -50.4080946438, -35.0078440092, -67.3261369391, 32.2106724154, 33.1026527036, 80.3973186259, 36.2330134377};
test_label[1623] = '{-67.3261369391};
test_output[1623] = '{147.723455565};
############ END DEBUG ############*/
test_input[12992:12999] = '{32'h41c77932, 32'hc2696338, 32'h426e017a, 32'hc287b9de, 32'h428e6cd9, 32'hc28c6aa0, 32'hc2a91ddb, 32'h4282a1ff};
test_label[1624] = '{32'hc287b9de};
test_output[1624] = '{32'h430b1410};
/*############ DEBUG ############
test_input[12992:12999] = '{24.9341771945, -58.3468939222, 59.5014423755, -67.8630217335, 71.2125966915, -70.208252629, -84.5583131538, 65.3163997479};
test_label[1624] = '{-67.8630217335};
test_output[1624] = '{139.078372713};
############ END DEBUG ############*/
test_input[13000:13007] = '{32'h4275180a, 32'h429cc135, 32'hc185133b, 32'h404e5b77, 32'hc0c2fb37, 32'hc2c6ce5a, 32'h42a63a2c, 32'hc24313ad};
test_label[1625] = '{32'hc24313ad};
test_output[1625] = '{32'h4303e43d};
/*############ DEBUG ############
test_input[13000:13007] = '{61.2734762048, 78.377354232, -16.6343894423, 3.22433253816, -6.09316608075, -99.4030274091, 83.1136152738, -48.7692134138};
test_label[1625] = '{-48.7692134138};
test_output[1625] = '{131.891561824};
############ END DEBUG ############*/
test_input[13008:13015] = '{32'h4277d765, 32'h41ff1fa3, 32'hc25d535b, 32'hc28fe2de, 32'h4295d884, 32'h42b57f7e, 32'h4200c8cd, 32'hc287afe9};
test_label[1626] = '{32'h4295d884};
test_output[1626] = '{32'h417d37cd};
/*############ DEBUG ############
test_input[13008:13015] = '{61.9603476356, 31.8904476174, -55.3314018619, -71.9430991193, 74.9228855673, 90.74900893, 32.1960956407, -67.8435750584};
test_label[1626] = '{74.9228855673};
test_output[1626] = '{15.8261234967};
############ END DEBUG ############*/
test_input[13016:13023] = '{32'h428fe71d, 32'hc2815705, 32'hc2aff7a7, 32'h4214704f, 32'h426fd833, 32'hc2433439, 32'h426c3f94, 32'hc28e56f3};
test_label[1627] = '{32'hc28e56f3};
test_output[1627] = '{32'h430f1f09};
/*############ DEBUG ############
test_input[13016:13023] = '{71.9513895459, -64.6699569723, -87.9836954875, 37.1096778332, 59.9611327281, -48.8009975242, 59.0620889658, -71.1698255651};
test_label[1627] = '{-71.1698255651};
test_output[1627] = '{143.12122384};
############ END DEBUG ############*/
test_input[13024:13031] = '{32'hc2a11c62, 32'hc2b56101, 32'hc1fb6ce0, 32'hc1d42db2, 32'h41d850f1, 32'h429d5526, 32'hc2a2caa1, 32'hc0d2ebec};
test_label[1628] = '{32'hc2a2caa1};
test_output[1628] = '{32'h43200fe3};
/*############ DEBUG ############
test_input[13024:13031] = '{-80.5554349494, -90.689461162, -31.4281622025, -26.5223128579, 27.0395229041, 78.6663057499, -81.3957570533, -6.59129929016};
test_label[1628] = '{-81.3957570533};
test_output[1628] = '{160.062062803};
############ END DEBUG ############*/
test_input[13032:13039] = '{32'hc1975742, 32'h4297d341, 32'h426e9754, 32'hc2689709, 32'hc1de994c, 32'hc147c6aa, 32'h420802cd, 32'h42849a1f};
test_label[1629] = '{32'h42849a1f};
test_output[1629] = '{32'h4119c956};
/*############ DEBUG ############
test_input[13032:13039] = '{-18.9176054542, 75.912607611, 59.6477815824, -58.1474966295, -27.8248517923, -12.4860015301, 34.002734206, 66.3010200629};
test_label[1629] = '{66.3010200629};
test_output[1629] = '{9.6116545807};
############ END DEBUG ############*/
test_input[13040:13047] = '{32'h4299ec05, 32'h42bdee9d, 32'h42171882, 32'h41fd168e, 32'h42221b64, 32'h416d3c6c, 32'hc23ab054, 32'hc201b210};
test_label[1630] = '{32'hc23ab054};
test_output[1630] = '{32'h430da363};
/*############ DEBUG ############
test_input[13040:13047] = '{76.9609749286, 94.9660411942, 37.773934188, 31.6360126318, 40.526749491, 14.8272517854, -46.6721937194, -32.4238877849};
test_label[1630] = '{-46.6721937194};
test_output[1630] = '{141.638234929};
############ END DEBUG ############*/
test_input[13048:13055] = '{32'h4189e3da, 32'h42a47472, 32'h408df481, 32'hc04c6004, 32'h425bac8d, 32'h42068c47, 32'hc183754b, 32'hc2389c3c};
test_label[1631] = '{32'h42068c47};
test_output[1631] = '{32'h42425c9d};
/*############ DEBUG ############
test_input[13048:13055] = '{17.2362549586, 82.2274323338, 4.43609671593, -3.19336036464, 54.9185059688, 33.6369895492, -16.4322724013, -46.1525718652};
test_label[1631] = '{33.6369895492};
test_output[1631] = '{48.5904427846};
############ END DEBUG ############*/
test_input[13056:13063] = '{32'hc2718093, 32'h42c17428, 32'hc2b65ed4, 32'h4131e398, 32'h420a7792, 32'h408d1a00, 32'h42afe6d9, 32'h425fa4b2};
test_label[1632] = '{32'h42afe6d9};
test_output[1632] = '{32'h410c6b1f};
/*############ DEBUG ############
test_input[13056:13063] = '{-60.3755604652, 96.7268709119, -91.1852092749, 11.1180649645, 34.6167694068, 4.4094237282, 87.9508730307, 55.910836572};
test_label[1632] = '{87.9508730307};
test_output[1632] = '{8.77615226412};
############ END DEBUG ############*/
test_input[13064:13071] = '{32'h420cf0d4, 32'h42bf1cd4, 32'hbe738054, 32'h41915d59, 32'hc208b5ee, 32'h4125f895, 32'h4217255d, 32'h416a318a};
test_label[1633] = '{32'h4125f895};
test_output[1633] = '{32'h42aa5dc1};
/*############ DEBUG ############
test_input[13064:13071] = '{35.2351818679, 95.5563028515, -0.237794225023, 18.1705803097, -34.177664707, 10.3731890369, 37.7864880877, 14.6370942946};
test_label[1633] = '{10.3731890369};
test_output[1633] = '{85.1831138146};
############ END DEBUG ############*/
test_input[13072:13079] = '{32'h42bd6609, 32'hc0c390cc, 32'hc0d31e84, 32'hc2ba9df3, 32'h42c5fc49, 32'h3f23b66b, 32'hc049af28, 32'h41089aad};
test_label[1634] = '{32'hc0d31e84};
test_output[1634] = '{32'h42d33523};
/*############ DEBUG ############
test_input[13072:13079] = '{94.6992876506, -6.11142544721, -6.5974751183, -93.3084924569, 98.9927406823, 0.639502208517, -3.15131576915, 8.53776284961};
test_label[1634] = '{-6.5974751183};
test_output[1634] = '{105.603781058};
############ END DEBUG ############*/
test_input[13080:13087] = '{32'hc14904a6, 32'h41c64458, 32'hc2951d40, 32'h4211c85a, 32'h426db07b, 32'h42a637d9, 32'h42762efd, 32'hc132098e};
test_label[1635] = '{32'hc14904a6};
test_output[1635] = '{32'h42bf586e};
/*############ DEBUG ############
test_input[13080:13087] = '{-12.5636353281, 24.7833713756, -74.5571296135, 36.4456549681, 59.4223456821, 83.1090785032, 61.5458869304, -11.1273331047};
test_label[1635] = '{-12.5636353281};
test_output[1635] = '{95.6727138318};
############ END DEBUG ############*/
test_input[13088:13095] = '{32'hc153cdd4, 32'h405ef823, 32'hc2867282, 32'h41aaaf2c, 32'h427156fb, 32'hc0f1f72e, 32'h427140ec, 32'hc28ba858};
test_label[1636] = '{32'hc2867282};
test_output[1636] = '{32'h43003db4};
/*############ DEBUG ############
test_input[13088:13095] = '{-13.2377508089, 3.48389499082, -67.2236466193, 21.3355325585, 60.3349433655, -7.56142337975, 60.3133993004, -69.8287992024};
test_label[1636] = '{-67.2236466193};
test_output[1636] = '{128.24102315};
############ END DEBUG ############*/
test_input[13096:13103] = '{32'hc29bc308, 32'h42ad6e95, 32'h40b22529, 32'h422e35f0, 32'hc265174e, 32'h421bd3ae, 32'h40b7d721, 32'h4294e814};
test_label[1637] = '{32'h421bd3ae};
test_output[1637] = '{32'h423f097e};
/*############ DEBUG ############
test_input[13096:13103] = '{-77.8809191832, 86.715982698, 5.56703622085, 43.5526747516, -57.2727579445, 38.9567171972, 5.74501061477, 74.4532742689};
test_label[1637] = '{38.9567171972};
test_output[1637] = '{47.7592702255};
############ END DEBUG ############*/
test_input[13104:13111] = '{32'hc2c050ee, 32'h426d0487, 32'h42020e3c, 32'hc2330685, 32'h4248aac5, 32'h4242c3b6, 32'h42b34adc, 32'h4296e043};
test_label[1638] = '{32'h4296e043};
test_output[1638] = '{32'h416354ca};
/*############ DEBUG ############
test_input[13104:13111] = '{-96.158062821, 59.2544204715, 32.513902497, -44.7563681086, 50.1667683961, 48.6911244967, 89.6462128073, 75.438012915};
test_label[1638] = '{75.438012915};
test_output[1638] = '{14.2082005675};
############ END DEBUG ############*/
test_input[13112:13119] = '{32'hc28f2281, 32'h42651b68, 32'hc24e0dd9, 32'hc2b2ae5f, 32'h40c207a4, 32'h4192faf1, 32'h426168d7, 32'hc26f87fd};
test_label[1639] = '{32'h4192faf1};
test_output[1639] = '{32'h421cf41f};
/*############ DEBUG ############
test_input[13112:13119] = '{-71.5673886939, 57.276762567, -51.5135242509, -89.3405660687, 6.06343272779, 18.3725304454, 56.352382052, -59.882801905};
test_label[1639] = '{18.3725304454};
test_output[1639] = '{39.238399662};
############ END DEBUG ############*/
test_input[13120:13127] = '{32'hc2a1fc57, 32'h42095b0f, 32'h42c75eda, 32'hc28828ef, 32'hc292c2b4, 32'h42ac617f, 32'hc2888624, 32'h4214a9af};
test_label[1640] = '{32'h4214a9af};
test_output[1640] = '{32'h427a1405};
/*############ DEBUG ############
test_input[13120:13127] = '{-80.9928488952, 34.3389240256, 99.6852569755, -68.0799456849, -73.3802777798, 86.1904184586, -68.2619903506, 37.1657072896};
test_label[1640] = '{37.1657072896};
test_output[1640] = '{62.5195510639};
############ END DEBUG ############*/
test_input[13128:13135] = '{32'h42bee5cc, 32'hc280921d, 32'hc15771d3, 32'hc24fa11e, 32'h4206c36f, 32'h421bd564, 32'hc2b448ff, 32'hc207c3bd};
test_label[1641] = '{32'hc24fa11e};
test_output[1641] = '{32'h43135b2d};
/*############ DEBUG ############
test_input[13128:13135] = '{95.4488203038, -64.2853743318, -13.4652891193, -51.907339933, 33.6908532462, 38.9583890389, -90.14256726, -33.9411518851};
test_label[1641] = '{-51.907339933};
test_output[1641] = '{147.356160237};
############ END DEBUG ############*/
test_input[13136:13143] = '{32'h42188bcd, 32'hc1916c8e, 32'h42c0e94e, 32'hc2a82bd1, 32'hc02df391, 32'hc18565ca, 32'h41299fef, 32'hc18d646f};
test_label[1642] = '{32'hc2a82bd1};
test_output[1642] = '{32'h43348a8f};
/*############ DEBUG ############
test_input[13136:13143] = '{38.13652405, -18.1780056324, 96.4556709187, -84.0855774213, -2.71799122203, -16.6747026144, 10.601546703, -17.6740399652};
test_label[1642] = '{-84.0855774213};
test_output[1642] = '{180.54124834};
############ END DEBUG ############*/
test_input[13144:13151] = '{32'hc1e38a12, 32'h40fb9653, 32'hc200c3fa, 32'h41dc4a0a, 32'h427d7b20, 32'h427c8dec, 32'h420333ef, 32'hc0fe7bfc};
test_label[1643] = '{32'h41dc4a0a};
test_output[1643] = '{32'h4211ac24};
/*############ DEBUG ############
test_input[13144:13151] = '{-28.4424179676, 7.86210027896, -32.1913838365, 27.5361523081, 63.3702380596, 63.1385966125, 32.8007177972, -7.9526347671};
test_label[1643] = '{27.5361523081};
test_output[1643] = '{36.4181044863};
############ END DEBUG ############*/
test_input[13152:13159] = '{32'h428d5dd5, 32'hc1c5c523, 32'h42942c3c, 32'h428917cf, 32'hc2ad74e1, 32'h429264f7, 32'h403eadc3, 32'hc0c6d0c2};
test_label[1644] = '{32'h428d5dd5};
test_output[1644] = '{32'h40718013};
/*############ DEBUG ############
test_input[13152:13159] = '{70.6832624007, -24.7212573127, 74.0863972355, 68.5464975862, -86.7282808854, 73.197195065, 2.97935560709, -6.21298336906};
test_label[1644] = '{70.6832624007};
test_output[1644] = '{3.77344191376};
############ END DEBUG ############*/
test_input[13160:13167] = '{32'hc23ca07e, 32'h4209e0f7, 32'h408f7dfc, 32'hc2486588, 32'h42a2d8b9, 32'h41bf7c46, 32'h42815bd5, 32'h4271da0e};
test_label[1645] = '{32'h42815bd5};
test_output[1645] = '{32'h4185f392};
/*############ DEBUG ############
test_input[13160:13167] = '{-47.1567324523, 34.4696939853, 4.48412881337, -50.0991512923, 81.4232901299, 23.9356812976, 64.679358948, 60.4629459007};
test_label[1645] = '{64.679358948};
test_output[1645] = '{16.7439312362};
############ END DEBUG ############*/
test_input[13168:13175] = '{32'h42077a12, 32'h417839c5, 32'h41a037b0, 32'h4166a3d3, 32'hc0268f3a, 32'hc2bead74, 32'hc198256e, 32'hc1c604e4};
test_label[1646] = '{32'hc0268f3a};
test_output[1646] = '{32'h4211e306};
/*############ DEBUG ############
test_input[13168:13175] = '{33.869209937, 15.5141042265, 20.0271913974, 14.4149959615, -2.60249197222, -95.3387760206, -19.0182768142, -24.7523884826};
test_label[1646] = '{-2.60249197222};
test_output[1646] = '{36.4717028973};
############ END DEBUG ############*/
test_input[13176:13183] = '{32'hc2bfca01, 32'hc2a930ff, 32'hc0477206, 32'hc1cc851a, 32'h421987ab, 32'hc102832c, 32'h41f8d071, 32'h41a4f4cb};
test_label[1647] = '{32'hc102832c};
test_output[1647] = '{32'h423a292b};
/*############ DEBUG ############
test_input[13176:13183] = '{-95.8945362696, -84.5956975747, -3.11633433924, -25.5649915167, 38.3824892778, -8.15702425781, 31.1017786314, 20.6195279421};
test_label[1647] = '{-8.15702425781};
test_output[1647] = '{46.5402020139};
############ END DEBUG ############*/
test_input[13184:13191] = '{32'h420ad096, 32'hc1ea7913, 32'hc1ca6949, 32'hc29c60cf, 32'hc0894be9, 32'hc1922a49, 32'hc2b7787e, 32'hc266c34c};
test_label[1648] = '{32'hc1922a49};
test_output[1648] = '{32'h4253e5bb};
/*############ DEBUG ############
test_input[13184:13191] = '{34.7036984559, -29.3091182134, -25.3014078157, -78.1890827196, -4.29051643156, -18.2706474452, -91.7353386694, -57.6907214234};
test_label[1648] = '{-18.2706474452};
test_output[1648] = '{52.974345901};
############ END DEBUG ############*/
test_input[13192:13199] = '{32'hc2bbd103, 32'h41e94434, 32'h42a9f145, 32'hc2335d97, 32'h426bada4, 32'h425c5b21, 32'hc1c8f64f, 32'hc16a3d4b};
test_label[1649] = '{32'h41e94434};
test_output[1649] = '{32'h425f4070};
/*############ DEBUG ############
test_input[13192:13199] = '{-93.9082242286, 29.1583019191, 84.9712295513, -44.8413965844, 58.9195714765, 55.088992861, -25.1202681828, -14.6399641929};
test_label[1649] = '{29.1583019191};
test_output[1649] = '{55.8129276322};
############ END DEBUG ############*/
test_input[13200:13207] = '{32'h428873bd, 32'hc21a9d71, 32'hc2061b3f, 32'hc2159e2f, 32'hc1eb587b, 32'hc2ab27fa, 32'h425b6358, 32'hc2a591db};
test_label[1650] = '{32'hc2159e2f};
test_output[1650] = '{32'h42d342d5};
/*############ DEBUG ############
test_input[13200:13207] = '{68.2260551363, -38.6537531355, -33.5266082077, -37.4044776709, -29.4182030753, -85.5780818525, 54.8470148919, -82.784872671};
test_label[1650] = '{-37.4044776709};
test_output[1650] = '{105.630534354};
############ END DEBUG ############*/
test_input[13208:13215] = '{32'hc2b36f6e, 32'hc178d879, 32'hc2ab10b2, 32'hc2aaa28f, 32'hc224444b, 32'h42347aef, 32'h42bd7cb6, 32'hc2562379};
test_label[1651] = '{32'h42bd7cb6};
test_output[1651] = '{32'h80000000};
/*############ DEBUG ############
test_input[13208:13215] = '{-89.7176365099, -15.5528497156, -85.5326108214, -85.3174994848, -41.0666907991, 45.1200537013, 94.7435730682, -53.5346397355};
test_label[1651] = '{94.7435730682};
test_output[1651] = '{-0.0};
############ END DEBUG ############*/
test_input[13216:13223] = '{32'hc17f23e3, 32'hc05eac02, 32'hc2a1774e, 32'hc2a7f155, 32'h42974ea6, 32'hc22308c5, 32'h42566cfe, 32'hc10446ff};
test_label[1652] = '{32'hc17f23e3};
test_output[1652] = '{32'h42b73323};
/*############ DEBUG ############
test_input[13216:13223] = '{-15.9462612386, -3.47924863009, -80.733014069, -83.9713503969, 75.6536116071, -40.7585634142, 53.606437752, -8.26733327731};
test_label[1652] = '{-15.9462612386};
test_output[1652] = '{91.5998728459};
############ END DEBUG ############*/
test_input[13224:13231] = '{32'hc2374e8a, 32'h421f8c8f, 32'h41a76d26, 32'hc1c383c7, 32'h42c1a2a9, 32'hc291699f, 32'hbfe8fede, 32'h4204e289};
test_label[1653] = '{32'h42c1a2a9};
test_output[1653] = '{32'h80000000};
/*############ DEBUG ############
test_input[13224:13231] = '{-45.8266989876, 39.8872644348, 20.9282943965, -24.4393444943, 96.8176956659, -72.7062887498, -1.82027795785, 33.2212250068};
test_label[1653] = '{96.8176956659};
test_output[1653] = '{-0.0};
############ END DEBUG ############*/
test_input[13232:13239] = '{32'h424d303b, 32'hc1e15cc1, 32'hc251d41b, 32'hc2311007, 32'hc21d3295, 32'hc27b7bba, 32'h4269169a, 32'h41a2229f};
test_label[1654] = '{32'hc21d3295};
test_output[1654] = '{32'h42c32512};
/*############ DEBUG ############
test_input[13232:13239] = '{51.2971018098, -28.1702893859, -52.4571327164, -44.2656531503, -39.2993966568, -62.8708273073, 58.2720713676, 20.2669042864};
test_label[1654] = '{-39.2993966568};
test_output[1654] = '{97.5724025823};
############ END DEBUG ############*/
test_input[13240:13247] = '{32'h427231e1, 32'h41e8b7b5, 32'h42681c3f, 32'hc28207d0, 32'h421805bc, 32'hc108d7d8, 32'hc23103c2, 32'h4228ef57};
test_label[1655] = '{32'h4228ef57};
test_output[1655] = '{32'h41932366};
/*############ DEBUG ############
test_input[13240:13247] = '{60.5487117335, 29.0896999207, 58.0275832019, -65.0152561075, 38.0056014123, -8.55269665397, -44.2536704676, 42.2337303304};
test_label[1655] = '{42.2337303304};
test_output[1655] = '{18.3922839304};
############ END DEBUG ############*/
test_input[13248:13255] = '{32'hc2867fc8, 32'hc18972c3, 32'h425de70e, 32'h421d61c2, 32'h423839b3, 32'h41c2d009, 32'hc2c3c33b, 32'h4276c5a6};
test_label[1656] = '{32'hc18972c3};
test_output[1656] = '{32'h429dc089};
/*############ DEBUG ############
test_input[13248:13255] = '{-67.2495728784, -17.1810362281, 55.4756383082, 39.3454673752, 46.0563465406, 24.3515804295, -97.8813102439, 61.6930179085};
test_label[1656] = '{-17.1810362281};
test_output[1656] = '{78.8760467767};
############ END DEBUG ############*/
test_input[13256:13263] = '{32'h42156245, 32'h426ba6bf, 32'h41b935b5, 32'h42c629a7, 32'hc287a53c, 32'h41cd7d18, 32'h42518e4f, 32'h41ba0daf};
test_label[1657] = '{32'h41b935b5};
test_output[1657] = '{32'h4297dc3a};
/*############ DEBUG ############
test_input[13256:13263] = '{37.3459665068, 58.9128383702, 23.1512249178, 99.0813516652, -67.8227200238, 25.6860800638, 52.3889732423, 23.2566804988};
test_label[1657] = '{23.1512249178};
test_output[1657] = '{75.9301267473};
############ END DEBUG ############*/
test_input[13264:13271] = '{32'hc2ab5c06, 32'hc237045e, 32'h42036438, 32'hc1d47dcb, 32'h3f86526f, 32'h420e2abe, 32'h42bb8913, 32'hc2a557dd};
test_label[1658] = '{32'h420e2abe};
test_output[1658] = '{32'h4268e769};
/*############ DEBUG ############
test_input[13264:13271] = '{-85.6797356374, -45.7542644685, 32.8478699931, -26.5614229008, 1.04939065442, 35.541739176, 93.767725058, -82.6716063298};
test_label[1658] = '{35.541739176};
test_output[1658] = '{58.225985882};
############ END DEBUG ############*/
test_input[13272:13279] = '{32'hc2517f54, 32'h4201bd0b, 32'hc20ffd1b, 32'h3fcf2f9a, 32'hc2a51b93, 32'h42bb40d0, 32'h40eaa3cd, 32'hc2b007b6};
test_label[1659] = '{32'hc2517f54};
test_output[1659] = '{32'h4312003d};
/*############ DEBUG ############
test_input[13272:13279] = '{-52.3743431488, 32.4346117413, -35.9971725413, 1.61864018379, -82.5538544361, 93.6265831662, 7.33249525633, -88.0150576153};
test_label[1659] = '{-52.3743431488};
test_output[1659] = '{146.000926315};
############ END DEBUG ############*/
test_input[13280:13287] = '{32'hc26d67d5, 32'h41c2b716, 32'hc1b2d22d, 32'h42a17d00, 32'h42ad98a6, 32'h41efff43, 32'hc2b96301, 32'h4283b777};
test_label[1660] = '{32'hc1b2d22d};
test_output[1660] = '{32'h42da4e64};
/*############ DEBUG ############
test_input[13280:13287] = '{-59.3513982723, 24.3393978986, -22.3526243305, 80.7441410116, 86.7981377131, 29.999639722, -92.693366307, 65.8583265687};
test_label[1660] = '{-22.3526243305};
test_output[1660] = '{109.153107748};
############ END DEBUG ############*/
test_input[13288:13295] = '{32'hc2931920, 32'hc001a7a6, 32'h4257f6dc, 32'hc296777f, 32'hc1fcfde7, 32'h42a0a9b9, 32'h42b06d8e, 32'hc1f6d857};
test_label[1661] = '{32'hc1f6d857};
test_output[1661] = '{32'h42ee23d5};
/*############ DEBUG ############
test_input[13288:13295] = '{-73.5490721471, -2.02585751075, 53.9910735752, -75.2333890823, -31.6239755282, 80.3314899861, 88.2139730681, -30.8556337651};
test_label[1661] = '{-30.8556337651};
test_output[1661] = '{119.069984057};
############ END DEBUG ############*/
test_input[13296:13303] = '{32'h421b12e5, 32'h426b5774, 32'hc292c7f3, 32'h429518f3, 32'hc28f7451, 32'h41f927f2, 32'hc2821664, 32'h42641b9c};
test_label[1662] = '{32'h429518f3};
test_output[1662] = '{32'h343b5484};
/*############ DEBUG ############
test_input[13296:13303] = '{38.7684531935, 58.8354049614, -73.3905262558, 74.5487320776, -71.7271775731, 31.1445053732, -65.0437313107, 57.0269617579};
test_label[1662] = '{74.5487320776};
test_output[1662] = '{1.74464781964e-07};
############ END DEBUG ############*/
test_input[13304:13311] = '{32'h4227a0c0, 32'h42c222f0, 32'hc1a34f42, 32'h421e329f, 32'hc29086e5, 32'h4296f03b, 32'h421efe29, 32'h429afdce};
test_label[1663] = '{32'h421e329f};
test_output[1663] = '{32'h42661340};
/*############ DEBUG ############
test_input[13304:13311] = '{41.9069814555, 97.0682337439, -20.4137009029, 39.5494337565, -72.2634647029, 75.4692001606, 39.7482016051, 77.4957122684};
test_label[1663] = '{39.5494337565};
test_output[1663] = '{57.518799991};
############ END DEBUG ############*/
test_input[13312:13319] = '{32'hc1d6d201, 32'hc2241f1a, 32'hc1a7d3ce, 32'hc2461319, 32'h42c256fd, 32'h422a3cd3, 32'hc2af0150, 32'h3f6417e5};
test_label[1664] = '{32'hc2461319};
test_output[1664] = '{32'h4312b045};
/*############ DEBUG ############
test_input[13312:13319] = '{-26.8525403054, -41.0303718982, -20.9784210429, -49.5186517497, 97.1698973027, 42.5593982051, -87.5025642051, 0.890989607519};
test_label[1664] = '{-49.5186517497};
test_output[1664] = '{146.688549052};
############ END DEBUG ############*/
test_input[13320:13327] = '{32'hc275d557, 32'h42af6405, 32'hc2865209, 32'h41a61364, 32'h425181c7, 32'hc2c21d97, 32'h4293866d, 32'h4210fd03};
test_label[1665] = '{32'hc275d557};
test_output[1665] = '{32'h43152758};
/*############ DEBUG ############
test_input[13320:13327] = '{-61.4583378573, 87.6953521556, -67.1602243879, 20.7594673452, 52.3767344849, -97.057795192, 73.7625517146, 36.2470835803};
test_label[1665] = '{-61.4583378573};
test_output[1665] = '{149.153690902};
############ END DEBUG ############*/
test_input[13328:13335] = '{32'h42134f31, 32'hc1a841d0, 32'h4237c8a5, 32'h4243c1ad, 32'hc2b28b97, 32'hc13fb771, 32'h42005032, 32'h423aa308};
test_label[1666] = '{32'h42005032};
test_output[1666] = '{32'h41880582};
/*############ DEBUG ############
test_input[13328:13335] = '{36.8273342613, -21.0321340807, 45.9459426479, 48.9391357, -89.2726344289, -11.9822856206, 32.0783146235, 46.659211004};
test_label[1666] = '{32.0783146235};
test_output[1666] = '{17.0026891244};
############ END DEBUG ############*/
test_input[13336:13343] = '{32'h41df1f98, 32'hc2ad8a05, 32'hc26eedd6, 32'hc196b213, 32'h41f4d08a, 32'hc19a0889, 32'hc2b16ea4, 32'h429cead6};
test_label[1667] = '{32'h41f4d08a};
test_output[1667] = '{32'h423f6d67};
/*############ DEBUG ############
test_input[13336:13343] = '{27.8904272557, -86.7695664291, -59.7322619965, -18.8369505686, 30.6018249507, -19.254167676, -88.7160972934, 78.4586625219};
test_label[1667] = '{30.6018249507};
test_output[1667] = '{47.8568375712};
############ END DEBUG ############*/
test_input[13344:13351] = '{32'h42c338ba, 32'h4198d5eb, 32'h42abaf90, 32'h4243a045, 32'h4217988f, 32'hc1ceecfb, 32'hc26eda71, 32'hc13e3b02};
test_label[1668] = '{32'h4243a045};
test_output[1668] = '{32'h4242d131};
/*############ DEBUG ############
test_input[13344:13351] = '{97.6107937635, 19.1044528323, 85.8428973442, 48.9065124047, 37.8989825299, -25.8657123808, -59.7133235334, -11.8894058345};
test_label[1668] = '{48.9065124047};
test_output[1668] = '{48.7042891082};
############ END DEBUG ############*/
test_input[13352:13359] = '{32'hc2c57110, 32'hc2c04236, 32'hc2b9ae42, 32'h42079f19, 32'hc2bb3d01, 32'hc26dc839, 32'h423d4dcc, 32'hc2b498f3};
test_label[1669] = '{32'hc2b498f3};
test_output[1669] = '{32'h43099fec};
/*############ DEBUG ############
test_input[13352:13359] = '{-98.7208237857, -96.1293199657, -92.8403487197, 33.9053679677, -93.6191446226, -59.4455292775, 47.3259719989, -90.2987279074};
test_label[1669] = '{-90.2987279074};
test_output[1669] = '{137.624701391};
############ END DEBUG ############*/
test_input[13360:13367] = '{32'h4252157a, 32'hc2bc068c, 32'h426dfe37, 32'h3fd0cfa9, 32'h42c178d2, 32'h40c527c3, 32'h422117a9, 32'h42906d1e};
test_label[1670] = '{32'h4252157a};
test_output[1670] = '{32'h4230dc29};
/*############ DEBUG ############
test_input[13360:13367] = '{52.5209744009, -94.0127896406, 59.4982576312, 1.63133733561, 96.7359761007, 6.16110383931, 40.2731059386, 72.213119712};
test_label[1670] = '{52.5209744009};
test_output[1670] = '{44.2150016998};
############ END DEBUG ############*/
test_input[13368:13375] = '{32'hc0e692f4, 32'hc2b568ff, 32'h41ad0c6b, 32'h426cf383, 32'h416a7c8a, 32'h41fd4cf7, 32'hc1f52308, 32'hc230c909};
test_label[1671] = '{32'hc0e692f4};
test_output[1671] = '{32'h4284e2f1};
/*############ DEBUG ############
test_input[13368:13375] = '{-7.20543884241, -90.7050741245, 21.6310639256, 59.237803993, 14.6554054598, 31.6625806706, -30.6421058854, -44.196321991};
test_label[1671] = '{-7.20543884241};
test_output[1671] = '{66.4432428354};
############ END DEBUG ############*/
test_input[13376:13383] = '{32'h41f2f924, 32'h415e694c, 32'h40d1376f, 32'h4251ee08, 32'h42863342, 32'hc28c407a, 32'h426e2afe, 32'hc2301271};
test_label[1672] = '{32'h42863342};
test_output[1672] = '{32'h3a08e1ae};
/*############ DEBUG ############
test_input[13376:13383] = '{30.3716515952, 13.9007067777, 6.53801688704, 52.4824531634, 67.1001147523, -70.1259324968, 59.5419838701, -44.0180091066};
test_label[1672] = '{67.1001147523};
test_output[1672] = '{0.000522161744836};
############ END DEBUG ############*/
test_input[13384:13391] = '{32'hc28a0979, 32'hc254841d, 32'h4293bb12, 32'h403aab14, 32'h41c64867, 32'hc298e35b, 32'hc1f4eccd, 32'h425c41c6};
test_label[1673] = '{32'h4293bb12};
test_output[1673] = '{32'h31eadd2a};
/*############ DEBUG ############
test_input[13384:13391] = '{-69.0185049832, -53.1290158407, 73.8653753144, 2.91669174405, 24.7853533052, -76.4440540245, -30.6156261012, 55.0642302863};
test_label[1673] = '{73.8653753144};
test_output[1673] = '{6.83543979312e-09};
############ END DEBUG ############*/
test_input[13392:13399] = '{32'hc127a547, 32'hc232960b, 32'h41ad2c18, 32'h42b5d6d8, 32'h412d4f3c, 32'hc206e2ad, 32'hc233504b, 32'hc2a5b235};
test_label[1674] = '{32'hc233504b};
test_output[1674] = '{32'h4307bf7f};
/*############ DEBUG ############
test_input[13392:13399] = '{-10.477850738, -44.6465263411, 21.6465297628, 90.9196144492, 10.8318443439, -33.7213614094, -44.8284110291, -82.8480573063};
test_label[1674] = '{-44.8284110291};
test_output[1674] = '{135.748025478};
############ END DEBUG ############*/
test_input[13400:13407] = '{32'h42255757, 32'hc28d010f, 32'h4118d6d2, 32'h42adac1f, 32'hc167c5c1, 32'h419aed97, 32'hc0b46bd7, 32'hc2900f46};
test_label[1675] = '{32'h42255757};
test_output[1675] = '{32'h423600e7};
/*############ DEBUG ############
test_input[13400:13407] = '{41.3352945955, -70.5020698725, 9.5524463044, 86.8361749395, -14.4857799247, 19.3660113249, -5.63816397383, -72.0298332366};
test_label[1675] = '{41.3352945955};
test_output[1675] = '{45.500880344};
############ END DEBUG ############*/
test_input[13408:13415] = '{32'h42b3af8a, 32'h4173b49d, 32'hc2140d62, 32'h416771fe, 32'hc29aa8f9, 32'h4296119b, 32'hc21e738e, 32'hc298c4d5};
test_label[1676] = '{32'hc29aa8f9};
test_output[1676] = '{32'h43272c42};
/*############ DEBUG ############
test_input[13408:13415] = '{89.8428533835, 15.2315946234, -37.0130698107, 14.4653304772, -77.3300225457, 75.0343868796, -39.612847789, -76.384437408};
test_label[1676] = '{-77.3300225457};
test_output[1676] = '{167.1728763};
############ END DEBUG ############*/
test_input[13416:13423] = '{32'h41cfe2c1, 32'h428a3967, 32'hc282ada0, 32'h422d0a6b, 32'h42948901, 32'hc2b92b29, 32'hc22801bc, 32'hc12d9565};
test_label[1677] = '{32'h42948901};
test_output[1677] = '{32'h3bbc7477};
/*############ DEBUG ############
test_input[13416:13423] = '{25.9857203008, 69.1121146465, -65.3391118458, 43.2601756102, 74.2675864451, -92.5842992123, -42.0016952431, -10.8489730405};
test_label[1677] = '{74.2675864451};
test_output[1677] = '{0.00575118837883};
############ END DEBUG ############*/
test_input[13424:13431] = '{32'h422b67f0, 32'h415de77e, 32'h3f41048d, 32'hc0b9513d, 32'hc220345e, 32'h41d92b56, 32'h42aef045, 32'h417f75ab};
test_label[1678] = '{32'h41d92b56};
test_output[1678] = '{32'h42714ade};
/*############ DEBUG ############
test_input[13424:13431] = '{42.8515004568, 13.8690166742, 0.753975686315, -5.79116679347, -40.0511382666, 27.1461604927, 87.4692733296, 15.9662273247};
test_label[1678] = '{27.1461604927};
test_output[1678] = '{60.323112837};
############ END DEBUG ############*/
test_input[13432:13439] = '{32'h425a0ebe, 32'hc244b4dd, 32'hc2b59557, 32'h4285fdc0, 32'hc2673e63, 32'hc28a1528, 32'hc28895f5, 32'hc1627304};
test_label[1679] = '{32'hc28895f5};
test_output[1679] = '{32'h430749db};
/*############ DEBUG ############
test_input[13432:13439] = '{54.5143949202, -49.1766256052, -90.7916784953, 66.9956082484, -57.8109233958, -69.0413212213, -68.2928879753, -14.1530804045};
test_label[1679] = '{-68.2928879753};
test_output[1679] = '{135.288500021};
############ END DEBUG ############*/
test_input[13440:13447] = '{32'h42481d90, 32'h42af60da, 32'h409f7a02, 32'h41da3370, 32'h425755bc, 32'h4108cf98, 32'hc203cf9b, 32'h42aa2b46};
test_label[1680] = '{32'h41da3370};
test_output[1680] = '{32'h4271f106};
/*############ DEBUG ############
test_input[13440:13447] = '{50.0288708439, 87.6891651725, 4.98364365913, 27.2751150711, 53.8337237506, 8.5506815942, -32.9527386692, 85.0845192197};
test_label[1680] = '{27.2751150711};
test_output[1680] = '{60.4853742732};
############ END DEBUG ############*/
test_input[13448:13455] = '{32'h41a2b17b, 32'hc2a20a55, 32'hc2c7c923, 32'hc1e2c94b, 32'hc22b554b, 32'hc216699d, 32'hc2ae22bd, 32'h40d06f68};
test_label[1681] = '{32'hc22b554b};
test_output[1681] = '{32'h427cae09};
/*############ DEBUG ############
test_input[13448:13455] = '{20.3366612109, -81.0201772213, -99.8928488949, -28.3482869625, -42.8332956827, -37.6031367002, -87.0678449884, 6.51359916836};
test_label[1681] = '{-42.8332956827};
test_output[1681] = '{63.1699578861};
############ END DEBUG ############*/
test_input[13456:13463] = '{32'h4299e18a, 32'hc28198f1, 32'h42bb8985, 32'h42a68e76, 32'hc24a6030, 32'h42c14930, 32'hc2a2da3b, 32'h4249384f};
test_label[1682] = '{32'h42bb8985};
test_output[1682] = '{32'h403b7929};
/*############ DEBUG ############
test_input[13456:13463] = '{76.9405058819, -64.798712033, 93.7685959509, 83.2782474873, -50.5939314186, 96.6429476315, -81.4262322115, 50.3049878998};
test_label[1682] = '{93.7685959509};
test_output[1682] = '{2.92926998111};
############ END DEBUG ############*/
test_input[13464:13471] = '{32'h42837610, 32'hc2a167fc, 32'h41b1739d, 32'h41d1ddec, 32'hc108d2a1, 32'hc2206789, 32'h42bd6422, 32'hc28265bc};
test_label[1683] = '{32'hc28265bc};
test_output[1683] = '{32'h431fe4ef};
/*############ DEBUG ############
test_input[13464:13471] = '{65.7305941039, -80.7030912371, 22.1814510806, 26.2333604941, -8.55142261755, -40.1011098705, 94.6955684839, -65.1986990912};
test_label[1683] = '{-65.1986990912};
test_output[1683] = '{159.894267575};
############ END DEBUG ############*/
test_input[13472:13479] = '{32'hc02b65c0, 32'h41dbe693, 32'h40c174ea, 32'h4282e3e6, 32'hc29515fa, 32'hc2bdc39d, 32'hc27b3896, 32'hc27ec35e};
test_label[1684] = '{32'h41dbe693};
test_output[1684] = '{32'h4217d482};
/*############ DEBUG ############
test_input[13472:13479] = '{-2.67808528676, 27.4875842409, 6.04552172037, 65.4451125825, -74.5429267285, -94.8820572151, -62.8052599293, -63.6907879724};
test_label[1684] = '{27.4875842409};
test_output[1684] = '{37.9575283416};
############ END DEBUG ############*/
test_input[13480:13487] = '{32'hc2c09dcb, 32'h427e399a, 32'hc218d790, 32'hc2c77ea2, 32'h414ab192, 32'h42c6c138, 32'h429c979c, 32'h428b099a};
test_label[1685] = '{32'hc2c09dcb};
test_output[1685] = '{32'h4343af81};
/*############ DEBUG ############
test_input[13480:13487] = '{-96.3081864421, 63.5562532456, -38.2105106329, -99.7473275227, 12.6683523133, 99.3773812078, 78.2961107015, 69.5187552842};
test_label[1685] = '{-96.3081864421};
test_output[1685] = '{195.685567651};
############ END DEBUG ############*/
test_input[13488:13495] = '{32'h42b0b131, 32'h4143bd6a, 32'h4146a4f7, 32'h42c3093d, 32'h4233b203, 32'h428051db, 32'h42bc1b95, 32'hc0ff0761};
test_label[1686] = '{32'h4233b203};
test_output[1686] = '{32'h42528021};
/*############ DEBUG ############
test_input[13488:13495] = '{88.3460751232, 12.2337432123, 12.4152747897, 97.5180454684, 44.9238388187, 64.1598743651, 94.0538738023, -7.96965064116};
test_label[1686] = '{44.9238388187};
test_output[1686] = '{52.6251264983};
############ END DEBUG ############*/
test_input[13496:13503] = '{32'hc29c3ef2, 32'hc264fa4c, 32'hc27970db, 32'h428c256b, 32'hc0e04798, 32'hc25c3e9e, 32'hc27852a8, 32'h42717161};
test_label[1687] = '{32'h428c256b};
test_output[1687] = '{32'h387de06f};
/*############ DEBUG ############
test_input[13496:13503] = '{-78.1229410496, -57.2444287909, -62.3602104654, 70.0730794786, -7.00873965345, -55.061150161, -62.0807197117, 60.360720448};
test_label[1687] = '{70.0730794786};
test_output[1687] = '{6.05289197168e-05};
############ END DEBUG ############*/
test_input[13504:13511] = '{32'h424828d4, 32'hc2a54ef5, 32'h4254de29, 32'h42bfd17d, 32'h403d6adb, 32'hc2a2e3ee, 32'h41f1bf0f, 32'h412180e5};
test_label[1688] = '{32'h412180e5};
test_output[1688] = '{32'h42aba161};
/*############ DEBUG ############
test_input[13504:13511] = '{50.0398722362, -82.6542157144, 53.2169519398, 95.9091583147, 2.95964689442, -81.445176522, 30.2182895926, 10.0939688245};
test_label[1688] = '{10.0939688245};
test_output[1688] = '{85.8151894902};
############ END DEBUG ############*/
test_input[13512:13519] = '{32'hc19927e0, 32'h422e25ab, 32'h42aff8fe, 32'hc1684c3b, 32'hc104fd58, 32'hc20c2edc, 32'hc2ac08b4, 32'h4122d8f4};
test_label[1689] = '{32'hc2ac08b4};
test_output[1689] = '{32'h432e00d9};
/*############ DEBUG ############
test_input[13512:13519] = '{-19.1444692941, 43.5367854599, 87.98630977, -14.5186111624, -8.31185172258, -35.0457626616, -86.0170000863, 10.1779666766};
test_label[1689] = '{-86.0170000863};
test_output[1689] = '{174.003309856};
############ END DEBUG ############*/
test_input[13520:13527] = '{32'h42c09a34, 32'h42736931, 32'hc27c56f9, 32'hc27889e6, 32'hc2589b39, 32'hc1cc477e, 32'hc2a8e9a7, 32'h4296faf0};
test_label[1690] = '{32'hc27c56f9};
test_output[1690] = '{32'h431f62d8};
/*############ DEBUG ############
test_input[13520:13527] = '{96.3011746663, 60.8527265097, -63.0849334915, -62.13466755, -54.1515838829, -25.5349074123, -84.4563560334, 75.4901099179};
test_label[1690] = '{-63.0849334915};
test_output[1690] = '{159.386108159};
############ END DEBUG ############*/
test_input[13528:13535] = '{32'h4064416e, 32'hc1f1c387, 32'h42499243, 32'hc2bf09ad, 32'h416cf247, 32'hc28ecfdf, 32'hc2b710f0, 32'hc2117cb2};
test_label[1691] = '{32'h4064416e};
test_output[1691] = '{32'h423b4e2c};
/*############ DEBUG ############
test_input[13528:13535] = '{3.56649341946, -30.2204713838, 50.3928346216, -95.5188962318, 14.8091500484, -71.4059952957, -91.5330828555, -36.3717725006};
test_label[1691] = '{3.56649341946};
test_output[1691] = '{46.8263412021};
############ END DEBUG ############*/
test_input[13536:13543] = '{32'hc251c62d, 32'hc2ac5e43, 32'h42b43ef6, 32'hc274cc0e, 32'h421515e7, 32'hc25feede, 32'hc18373e6, 32'hc117cd81};
test_label[1692] = '{32'hc251c62d};
test_output[1692] = '{32'h430e9107};
/*############ DEBUG ############
test_input[13536:13543] = '{-52.4435321387, -86.1841034933, 90.1229734126, -61.1992711414, 37.2713904996, -55.9832672404, -16.4315905702, -9.48767219753};
test_label[1692] = '{-52.4435321387};
test_output[1692] = '{142.566505551};
############ END DEBUG ############*/
test_input[13544:13551] = '{32'hc2a02c03, 32'h425aa76b, 32'h4283a64c, 32'hc18f9d93, 32'hc2aaf3d8, 32'hc17de8ef, 32'hc2152477, 32'h42a75e71};
test_label[1693] = '{32'hc2a02c03};
test_output[1693] = '{32'h4323c53a};
/*############ DEBUG ############
test_input[13544:13551] = '{-80.0859591962, 54.6634936648, 65.824795191, -17.9519407939, -85.4762542596, -15.8693682304, -37.2856101047, 83.684455381};
test_label[1693] = '{-80.0859591962};
test_output[1693] = '{163.770414595};
############ END DEBUG ############*/
test_input[13552:13559] = '{32'h4033bdde, 32'hc29d4640, 32'hc2596f35, 32'hc2674f6e, 32'hc2829434, 32'hc1abfae4, 32'hc1b97959, 32'hc1d183eb};
test_label[1694] = '{32'hc2596f35};
test_output[1694] = '{32'h4264ab13};
/*############ DEBUG ############
test_input[13552:13559] = '{2.80846352156, -78.6372078401, -54.3586006323, -57.8275669788, -65.2894570052, -21.4975057806, -23.1842522358, -26.1894135761};
test_label[1694] = '{-54.3586006323};
test_output[1694] = '{57.1670641539};
############ END DEBUG ############*/
test_input[13560:13567] = '{32'h41c32fc6, 32'h42c1b7f8, 32'hc23fc5cc, 32'h4293205f, 32'hbd9cec65, 32'hc2b82caf, 32'hc2984fb6, 32'h41db7f86};
test_label[1695] = '{32'h42c1b7f8};
test_output[1695] = '{32'h2ea7d440};
/*############ DEBUG ############
test_input[13560:13567] = '{24.3983263794, 96.8593157056, -47.9431621742, 73.5632277673, -0.0766227593303, -92.0872763399, -76.1556889235, 27.4372682282};
test_label[1695] = '{96.8593157056};
test_output[1695] = '{7.63198393401e-11};
############ END DEBUG ############*/
test_input[13568:13575] = '{32'h41d4f478, 32'hc26170eb, 32'hc1709a2a, 32'h425b4964, 32'h42331e87, 32'h41e74481, 32'h429dbd47, 32'h414a150f};
test_label[1696] = '{32'hc26170eb};
test_output[1696] = '{32'h43073ade};
/*############ DEBUG ############
test_input[13568:13575] = '{26.6193699537, -56.3602728648, -15.037638102, 54.8216718693, 44.7798128378, 28.9084499965, 78.8696801383, 12.6301408707};
test_label[1696] = '{-56.3602728648};
test_output[1696] = '{135.229953003};
############ END DEBUG ############*/
test_input[13576:13583] = '{32'h42c088fd, 32'hc277a1ea, 32'h41bfc9d0, 32'h422850a3, 32'h4278f843, 32'hc226043a, 32'hc2a5c443, 32'hc26163ff};
test_label[1697] = '{32'hc2a5c443};
test_output[1697] = '{32'h433326a0};
/*############ DEBUG ############
test_input[13576:13583] = '{96.2675558658, -61.9081205522, 23.9735405854, 42.0787480197, 62.2424421059, -41.5041257562, -82.8833236622, -56.3476539664};
test_label[1697] = '{-82.8833236622};
test_output[1697] = '{179.150879528};
############ END DEBUG ############*/
test_input[13584:13591] = '{32'hc0ca223c, 32'hc1d6868a, 32'h41a72740, 32'h42b3a114, 32'h42b9c2c2, 32'h4291303d, 32'hc1a855ef, 32'hc2373a6c};
test_label[1698] = '{32'h41a72740};
test_output[1698] = '{32'h42901046};
/*############ DEBUG ############
test_input[13584:13591] = '{-6.31667911799, -26.8156921745, 20.8941640903, 89.814609287, 92.8803851683, 72.5942130849, -21.0419604536, -45.8070512461};
test_label[1698] = '{20.8941640903};
test_output[1698] = '{72.0317847661};
############ END DEBUG ############*/
test_input[13592:13599] = '{32'h42c31be8, 32'hc28f0be5, 32'h41501a78, 32'h42a75e62, 32'hbffc752f, 32'h41b89619, 32'hc26a7f1f, 32'hc2881844};
test_label[1699] = '{32'h41b89619};
test_output[1699] = '{32'h4294f662};
/*############ DEBUG ############
test_input[13592:13599] = '{97.5545079544, -71.5232279455, 13.0064619214, 83.6843404804, -1.97232613721, 23.073289789, -58.6241405998, -68.0473959859};
test_label[1699] = '{23.073289789};
test_output[1699] = '{74.4812191122};
############ END DEBUG ############*/
test_input[13600:13607] = '{32'h4140c1cf, 32'hc29b3d08, 32'hc1c7f3d6, 32'hc2988b93, 32'h4142be3c, 32'hc2978214, 32'hc23c282d, 32'h423cd2b9};
test_label[1700] = '{32'hc2978214};
test_output[1700] = '{32'h42f5eb71};
/*############ DEBUG ############
test_input[13600:13607] = '{12.0473166279, -77.6191981513, -24.9940598702, -76.2726057744, 12.1714436326, -75.7540624915, -47.0392326005, 47.2057826334};
test_label[1700] = '{-75.7540624915};
test_output[1700] = '{122.959845125};
############ END DEBUG ############*/
test_input[13608:13615] = '{32'hc238cc25, 32'hc0e75d0e, 32'h413ba2f5, 32'hc25d43d0, 32'h42514c39, 32'hc223098b, 32'hc24f5239, 32'hc0a19780};
test_label[1701] = '{32'hc223098b};
test_output[1701] = '{32'h42ba2ae2};
/*############ DEBUG ############
test_input[13608:13615] = '{-46.1993597678, -7.23010897713, 11.7272846471, -55.3162220134, 52.3244362491, -40.7593191636, -51.8302948659, -5.04974356858};
test_label[1701] = '{-40.7593191636};
test_output[1701] = '{93.0837554127};
############ END DEBUG ############*/
test_input[13616:13623] = '{32'hbf869f6b, 32'h428e98d5, 32'h40176927, 32'h421a3659, 32'h42a88707, 32'h42838963, 32'h427577ed, 32'h42c64208};
test_label[1702] = '{32'h42c64208};
test_output[1702] = '{32'h34bbec3c};
/*############ DEBUG ############
test_input[13616:13623] = '{-1.05174007253, 71.2984963617, 2.36579309127, 38.5530755605, 84.2637285782, 65.7683316425, 61.3671142695, 99.1289678228};
test_label[1702] = '{99.1289678228};
test_output[1702] = '{3.50033465967e-07};
############ END DEBUG ############*/
test_input[13624:13631] = '{32'hc0adcb4d, 32'hc190d942, 32'hc23c37a4, 32'hc26a1ce5, 32'h41f8ca28, 32'hc2bc2356, 32'h4187d241, 32'hc263c8dc};
test_label[1703] = '{32'hc0adcb4d};
test_output[1703] = '{32'h42121e7e};
/*############ DEBUG ############
test_input[13624:13631] = '{-5.43106715567, -18.1060836374, -47.0543383902, -58.5282183149, 31.0987082777, -94.0690169018, 16.9776623665, -56.9461517101};
test_label[1703] = '{-5.43106715567};
test_output[1703] = '{36.5297761701};
############ END DEBUG ############*/
test_input[13632:13639] = '{32'h42865e8e, 32'hc1dfbf58, 32'h4287bfe1, 32'h4215d154, 32'h4226b8c9, 32'hc2936920, 32'h4201316c, 32'hc15a42f8};
test_label[1704] = '{32'h4215d154};
test_output[1704] = '{32'h41f69d57};
/*############ DEBUG ############
test_input[13632:13639] = '{67.1846741352, -27.9684300281, 67.8747613428, 37.4544206321, 41.6804558697, -73.7053215382, 32.2982649805, -13.6413494161};
test_label[1704] = '{37.4544206321};
test_output[1704] = '{30.8268268505};
############ END DEBUG ############*/
test_input[13640:13647] = '{32'hc1b6bf8c, 32'h42adc49d, 32'h42089bca, 32'hc2a0aec6, 32'h42bb2edc, 32'h4175abcf, 32'hc1b2ae23, 32'h4259053b};
test_label[1705] = '{32'hc2a0aec6};
test_output[1705] = '{32'h432def21};
/*############ DEBUG ############
test_input[13640:13647] = '{-22.8435279867, 86.8840117052, 34.152137101, -80.3413508162, 93.5915205127, 15.3544454983, -22.3350275471, 54.2551084072};
test_label[1705] = '{-80.3413508162};
test_output[1705] = '{173.934092287};
############ END DEBUG ############*/
test_input[13648:13655] = '{32'hc21e1324, 32'h40bb41f1, 32'h411a5ecf, 32'h426206fa, 32'h41c24b42, 32'h429daa75, 32'h42790cd6, 32'h4283a4ff};
test_label[1706] = '{32'h429daa75};
test_output[1706] = '{32'h361a5c67};
/*############ DEBUG ############
test_input[13648:13655] = '{-39.5186902591, 5.85179931873, 9.64814645202, 56.5068123895, 24.2867473291, 78.8329263371, 62.2625337925, 65.8222573342};
test_label[1706] = '{78.8329263371};
test_output[1706] = '{2.30015733741e-06};
############ END DEBUG ############*/
test_input[13656:13663] = '{32'h418bdd8d, 32'hc241c868, 32'hc21f3f9f, 32'hc298e61a, 32'h4209688f, 32'hc1a00f19, 32'h428326ff, 32'hc2007e29};
test_label[1707] = '{32'hc21f3f9f};
test_output[1707] = '{32'h42d2c6ce};
/*############ DEBUG ############
test_input[13656:13663] = '{17.4831795534, -48.4457082535, -39.8121311757, -76.4494142255, 34.352109184, -20.0073724606, 65.5761629787, -32.1232023549};
test_label[1707] = '{-39.8121311757};
test_output[1707] = '{105.388294154};
############ END DEBUG ############*/
test_input[13664:13671] = '{32'hc159e8ed, 32'h4219a30f, 32'hc1db250e, 32'h4207a448, 32'hc24b71e5, 32'h40aec399, 32'hc27b0620, 32'hc08e1952};
test_label[1708] = '{32'hc24b71e5};
test_output[1708] = '{32'h42b29024};
/*############ DEBUG ############
test_input[13664:13671] = '{-13.6193669354, 38.4092365992, -27.3930935672, 33.9104302159, -50.8612267963, 5.46137667196, -62.755979587, -4.44059071214};
test_label[1708] = '{-50.8612267963};
test_output[1708] = '{89.2815242622};
############ END DEBUG ############*/
test_input[13672:13679] = '{32'hc26a2c0d, 32'h42afcd73, 32'hc1adebb9, 32'h42aa54b5, 32'hc1a9d8f7, 32'hc29b2d72, 32'hc28e50e9, 32'h418e6e89};
test_label[1709] = '{32'h418e6e89};
test_output[1709] = '{32'h428c51fb};
/*############ DEBUG ############
test_input[13672:13679] = '{-58.5430196403, 87.9012660217, -21.7400985436, 85.1654444007, -21.2309399102, -77.588763521, -71.1580246165, 17.8039713841};
test_label[1709] = '{17.8039713841};
test_output[1709] = '{70.1601198582};
############ END DEBUG ############*/
test_input[13680:13687] = '{32'h3f08c45c, 32'h41ff4338, 32'h41d70857, 32'hc123fdfb, 32'h42a42ab6, 32'h42147c92, 32'h424e664e, 32'h42b8f812};
test_label[1710] = '{32'h42b8f812};
test_output[1710] = '{32'h37ff0101};
/*############ DEBUG ############
test_input[13680:13687] = '{0.534246196954, 31.9078223386, 26.8790728433, -10.2495072041, 82.0834210277, 37.1216491847, 51.5999064032, 92.4845120618};
test_label[1710] = '{92.4845120618};
test_output[1710] = '{3.03988361899e-05};
############ END DEBUG ############*/
test_input[13688:13695] = '{32'hc223c222, 32'h4247dee9, 32'hc240fd0a, 32'hc1a007e6, 32'hc1b84e80, 32'h4292679f, 32'hc295adb4, 32'hc2646233};
test_label[1711] = '{32'hc2646233};
test_output[1711] = '{32'h43024c5c};
/*############ DEBUG ############
test_input[13688:13695] = '{-40.9395820471, 49.9676852762, -48.2471073954, -20.0038574596, -23.0383294976, 73.2023857295, -74.8392607805, -57.0958959675};
test_label[1711] = '{-57.0958959675};
test_output[1711] = '{130.298281697};
############ END DEBUG ############*/
test_input[13696:13703] = '{32'hc2ac3e67, 32'hc20fb812, 32'hc1c5a292, 32'h41db3f0d, 32'h428d804f, 32'h414ba05c, 32'hc17036e7, 32'h429f203f};
test_label[1712] = '{32'h414ba05c};
test_output[1712] = '{32'h4285ac47};
/*############ DEBUG ############
test_input[13696:13703] = '{-86.1218763963, -35.9297556647, -24.7043791862, 27.4057858761, 70.7506035275, 12.7266500831, -15.013403922, 79.5629805487};
test_label[1712] = '{12.7266500831};
test_output[1712] = '{66.8364793335};
############ END DEBUG ############*/
test_input[13704:13711] = '{32'h42910bd4, 32'hc22f6d62, 32'h41811d32, 32'h42738043, 32'hc213bdc6, 32'hc149878e, 32'hc228bfbe, 32'hc23139a3};
test_label[1713] = '{32'h42910bd4};
test_output[1713] = '{32'h37129883};
/*############ DEBUG ############
test_input[13704:13711] = '{72.523104094, -43.8568173733, 16.1392550048, 60.8752549141, -36.9353262453, -12.595594151, -42.1872477154, -44.3062869922};
test_label[1713] = '{72.523104094};
test_output[1713] = '{8.73778748201e-06};
############ END DEBUG ############*/
test_input[13712:13719] = '{32'h42bb3173, 32'h42a5c31a, 32'h41093ccc, 32'h42a05276, 32'h428bdd40, 32'h4171a933, 32'hc265aff8, 32'h42bdfdaa};
test_label[1714] = '{32'h42bdfdaa};
test_output[1714] = '{32'h3e61f1b3};
/*############ DEBUG ############
test_input[13712:13719] = '{93.5965783992, 82.8810554698, 8.57734276253, 80.1610588421, 69.932126447, 15.1038084519, -57.421844809, 94.9954340466};
test_label[1714] = '{94.9954340466};
test_output[1714] = '{0.220648569848};
############ END DEBUG ############*/
test_input[13720:13727] = '{32'h42b315c4, 32'h413389d9, 32'h42700a9a, 32'h40924ccd, 32'hc24b8b0f, 32'h41b3bca7, 32'h41a6f95b, 32'hc2c4c98e};
test_label[1715] = '{32'h41b3bca7};
test_output[1715] = '{32'h4286269a};
/*############ DEBUG ############
test_input[13720:13727] = '{89.5425105631, 11.2211545022, 60.0103533408, 4.57187530302, -50.8857978186, 22.4671154789, 20.8717547545, -98.3936605296};
test_label[1715] = '{22.4671154789};
test_output[1715] = '{67.0753950841};
############ END DEBUG ############*/
test_input[13728:13735] = '{32'h4036a2bd, 32'h41f7889a, 32'hc29ac701, 32'h418c9f15, 32'h3f9d0543, 32'hc005feb1, 32'h42b2740d, 32'h40e0c5f4};
test_label[1716] = '{32'h418c9f15};
test_output[1716] = '{32'h428f4c47};
/*############ DEBUG ############
test_input[13728:13735] = '{2.85368275718, 30.9416999978, -77.3886824329, 17.5776767794, 1.22672304614, -2.09367012514, 89.2266583422, 7.02416414179};
test_label[1716] = '{17.5776767794};
test_output[1716] = '{71.6489815628};
############ END DEBUG ############*/
test_input[13736:13743] = '{32'hc10daf28, 32'h4218c4d4, 32'hc2b13cd1, 32'hc24689ac, 32'hc2a9a416, 32'h4284a80f, 32'h42bc7a2f, 32'h429725b3};
test_label[1717] = '{32'hc2b13cd1};
test_output[1717] = '{32'h4336db80};
/*############ DEBUG ############
test_input[13736:13743] = '{-8.85526285803, 38.192215234, -88.618783916, -49.6344441044, -84.8204833446, 66.3282430414, 94.2386435806, 75.5736314224};
test_label[1717] = '{-88.618783916};
test_output[1717] = '{182.857427504};
############ END DEBUG ############*/
test_input[13744:13751] = '{32'hc22ba3c4, 32'hc29dde7a, 32'h42aa4eeb, 32'h42830502, 32'h41a49ed6, 32'h41fcffbb, 32'hc0410af3, 32'h428c0253};
test_label[1718] = '{32'hc22ba3c4};
test_output[1718] = '{32'h43001066};
/*############ DEBUG ############
test_input[13744:13751] = '{-42.9099261013, -78.934527191, 85.1541374775, 65.5097824628, 20.57755652, 31.624868108, -3.01629334315, 70.0045429293};
test_label[1718] = '{-42.9099261013};
test_output[1718] = '{128.064063845};
############ END DEBUG ############*/
test_input[13752:13759] = '{32'h420602d4, 32'hc2a6be33, 32'hc1ee31d2, 32'hc2a657ff, 32'hc19e9543, 32'hc2b74217, 32'h42b79ecb, 32'hc2863ff7};
test_label[1719] = '{32'hc2b74217};
test_output[1719] = '{32'h43377071};
/*############ DEBUG ############
test_input[13752:13759] = '{33.5027611066, -83.3714791372, -29.7743258695, -83.1718655741, -19.8228819746, -91.6290800558, 91.8101387086, -67.1249304447};
test_label[1719] = '{-91.6290800558};
test_output[1719] = '{183.439218764};
############ END DEBUG ############*/
test_input[13760:13767] = '{32'hc1217b47, 32'hc26b8294, 32'hc271ed13, 32'h42c303a2, 32'h41fb2480, 32'h4009838e, 32'h427326b4, 32'hc2512a2b};
test_label[1720] = '{32'hc271ed13};
test_output[1720] = '{32'h431dfd16};
/*############ DEBUG ############
test_input[13760:13767] = '{-10.0925970778, -58.8775172063, -60.4815192686, 97.5070943338, 31.3928225551, 2.14865440393, 60.7877944766, -52.2911787881};
test_label[1720] = '{-60.4815192686};
test_output[1720] = '{157.988613602};
############ END DEBUG ############*/
test_input[13768:13775] = '{32'hc22b2fc6, 32'hc23861b0, 32'hc1974090, 32'h4232b3c5, 32'h423eeeaa, 32'h4284f6b2, 32'h41d3bf71, 32'hc2aff37a};
test_label[1721] = '{32'hc1974090};
test_output[1721] = '{32'h42aac6d6};
/*############ DEBUG ############
test_input[13768:13775] = '{-42.7966537118, -46.0953985589, -18.9065245206, 44.6755566592, 47.7330701638, 66.4818305245, 26.4684779446, -87.9755386428};
test_label[1721] = '{-18.9065245206};
test_output[1721] = '{85.3883550527};
############ END DEBUG ############*/
test_input[13776:13783] = '{32'hc28a8bd9, 32'h42c74c86, 32'h42268d56, 32'h41862b53, 32'h428a94af, 32'h3f775239, 32'hc1fdd316, 32'h42833aad};
test_label[1722] = '{32'h42c74c86};
test_output[1722] = '{32'h2996c000};
/*############ DEBUG ############
test_input[13776:13783] = '{-69.2731409688, 99.6494628884, 41.6380231926, 16.7711544677, 69.290397504, 0.966098368243, -31.7280694718, 65.614603223};
test_label[1722] = '{99.6494628884};
test_output[1722] = '{6.69464483849e-14};
############ END DEBUG ############*/
test_input[13784:13791] = '{32'hc20fe97a, 32'hc2615663, 32'hc2a5d5df, 32'hc00535bc, 32'h40e97bad, 32'hc1b8d528, 32'hc286c047, 32'hc1eb50d1};
test_label[1723] = '{32'hc1b8d528};
test_output[1723] = '{32'h41f33440};
/*############ DEBUG ############
test_input[13784:13791] = '{-35.9780031842, -56.3343610079, -82.9177166909, -2.08140474639, 7.29634735559, -23.1040801442, -67.3755442101, -29.4144606204};
test_label[1723] = '{-23.1040801442};
test_output[1723] = '{30.4005120814};
############ END DEBUG ############*/
test_input[13792:13799] = '{32'hc05af3b0, 32'h42a541e7, 32'h42c01131, 32'hc0fb405a, 32'h42059ccb, 32'hc096fba2, 32'hc243ace0, 32'hc2817dfc};
test_label[1724] = '{32'hc096fba2};
test_output[1724] = '{32'h42c980ec};
/*############ DEBUG ############
test_input[13792:13799] = '{-3.42112341432, 82.6287162747, 96.0335784726, -7.85160543648, 33.4031169142, -4.71821698584, -48.9188236253, -64.7460652361};
test_label[1724] = '{-4.71821698584};
test_output[1724] = '{100.751796966};
############ END DEBUG ############*/
test_input[13800:13807] = '{32'h429b2abc, 32'hc2b0dfcc, 32'h428c017d, 32'h429fa8e0, 32'h42c22b62, 32'hc2aa4e36, 32'hc1b59bf3, 32'hc2b1ad00};
test_label[1725] = '{32'hc2b1ad00};
test_output[1725] = '{32'h4339ec31};
/*############ DEBUG ############
test_input[13800:13807] = '{77.5834627732, -88.4371037119, 70.0029047282, 79.8298327047, 97.0847287242, -85.1527581292, -22.7011467927, -88.8378902885};
test_label[1725] = '{-88.8378902885};
test_output[1725] = '{185.922619048};
############ END DEBUG ############*/
test_input[13808:13815] = '{32'hc174d7b1, 32'h41679341, 32'h41f44ef1, 32'h4135b375, 32'h42ac8674, 32'hc2bafe71, 32'hc16a4501, 32'hc29863ca};
test_label[1726] = '{32'h4135b375};
test_output[1726] = '{32'h4295d005};
/*############ DEBUG ############
test_input[13808:13815] = '{-15.3026593207, 14.4734509465, 30.5385453513, 11.3563128859, 86.2626028811, -93.4969528142, -14.6418466396, -76.1949029617};
test_label[1726] = '{11.3563128859};
test_output[1726] = '{74.9062899952};
############ END DEBUG ############*/
test_input[13816:13823] = '{32'hc28358c4, 32'h40598f81, 32'h425ceeea, 32'hc26e041a, 32'h408d76f3, 32'hc2af98e6, 32'h429448c1, 32'h42649f01};
test_label[1727] = '{32'hc28358c4};
test_output[1727] = '{32'h430bd0c3};
/*############ DEBUG ############
test_input[13816:13823] = '{-65.6733729695, 3.39938369337, 55.2333147649, -59.5040048503, 4.42077011372, -87.7986270213, 74.1420985181, 57.1552788188};
test_label[1727] = '{-65.6733729695};
test_output[1727] = '{139.815471536};
############ END DEBUG ############*/
test_input[13824:13831] = '{32'h42360e92, 32'hc237562d, 32'hc2bd8109, 32'h41d05ba4, 32'h41df2bea, 32'hc20b3df2, 32'hc231bba4, 32'hc0cc5214};
test_label[1728] = '{32'hc237562d};
test_output[1728] = '{32'h42b6b260};
/*############ DEBUG ############
test_input[13824:13831] = '{45.5142295392, -45.834155421, -94.7520241655, 26.0447469224, 27.8964425764, -34.8104925593, -44.4332436657, -6.3850192111};
test_label[1728] = '{-45.834155421};
test_output[1728] = '{91.348384986};
############ END DEBUG ############*/
test_input[13832:13839] = '{32'h4036731e, 32'h40830ff7, 32'h41de62ae, 32'h422c33f5, 32'h4290afbf, 32'hbf908f79, 32'hc24a77e0, 32'h426a8eee};
test_label[1729] = '{32'h41de62ae};
test_output[1729] = '{32'h42322e27};
/*############ DEBUG ############
test_input[13832:13839] = '{2.85077630684, 4.09569873654, 27.7981825208, 43.050740083, 72.3432506386, -1.12937845072, -50.6170670492, 58.6395779126};
test_label[1729] = '{27.7981825208};
test_output[1729] = '{44.5450692361};
############ END DEBUG ############*/
test_input[13840:13847] = '{32'hc25f0422, 32'h41e2d291, 32'h420956e7, 32'h42a6786c, 32'h3f821d16, 32'h427c8b13, 32'hc2ae41e0, 32'hc2c39bc5};
test_label[1730] = '{32'hc25f0422};
test_output[1730] = '{32'h430afd3e};
/*############ DEBUG ############
test_input[13840:13847] = '{-55.7540351752, 28.3528163953, 34.3348647364, 83.2351966206, 1.01651259202, 63.135815872, -87.1286589986, -97.8042363697};
test_label[1730] = '{-55.7540351752};
test_output[1730] = '{138.989231798};
############ END DEBUG ############*/
test_input[13848:13855] = '{32'h4267377c, 32'hc2213861, 32'hc2990710, 32'hc1d71497, 32'hc29d6139, 32'h411423a4, 32'hc0b69cca, 32'hc2a92c4a};
test_label[1731] = '{32'hc2a92c4a};
test_output[1731] = '{32'h430e6404};
/*############ DEBUG ############
test_input[13848:13855] = '{57.8041834876, -40.3050559635, -76.5137971404, -26.8850527659, -78.6898915488, 9.25870179808, -5.70663915614, -84.5865022144};
test_label[1731] = '{-84.5865022144};
test_output[1731] = '{142.390685702};
############ END DEBUG ############*/
test_input[13856:13863] = '{32'h408551ce, 32'h422dd239, 32'hc14fd562, 32'h40994008, 32'hc2c61d94, 32'h42bbf98c, 32'hc2abf0d3, 32'hc223920f};
test_label[1732] = '{32'hc2abf0d3};
test_output[1732] = '{32'h4333f52f};
/*############ DEBUG ############
test_input[13856:13863] = '{4.16623591283, 43.4552948487, -12.9895955657, 4.78906653938, -99.057773367, 93.9873944359, -85.9703581011, -40.8926359335};
test_label[1732] = '{-85.9703581011};
test_output[1732] = '{179.957752537};
############ END DEBUG ############*/
test_input[13864:13871] = '{32'hc29cd260, 32'hc2a9cb58, 32'h41cc8467, 32'h4229ee0e, 32'h41bc0a85, 32'h4269d466, 32'h429bc14f, 32'h427a1f9b};
test_label[1733] = '{32'h4229ee0e};
test_output[1733] = '{32'h420d9490};
/*############ DEBUG ############
test_input[13864:13871] = '{-78.4108870059, -84.897152378, 25.5646494125, 42.4824765729, 23.5051369914, 58.4574188431, 77.8775554905, 62.5308631904};
test_label[1733] = '{42.4824765729};
test_output[1733] = '{35.3950791376};
############ END DEBUG ############*/
test_input[13872:13879] = '{32'hc281dedb, 32'hc27671a1, 32'hc2c5b7df, 32'h42772cd8, 32'hc2b5bd63, 32'hc202d459, 32'h41de58d0, 32'h41395538};
test_label[1734] = '{32'h41395538};
test_output[1734] = '{32'h4248d78a};
/*############ DEBUG ############
test_input[13872:13879] = '{-64.9352669225, -61.6109642133, -98.8591208634, 61.793791666, -90.8698944543, -32.7073706566, 27.7933655606, 11.5833054866};
test_label[1734] = '{11.5833054866};
test_output[1734] = '{50.2104861794};
############ END DEBUG ############*/
test_input[13880:13887] = '{32'h42be8cda, 32'h428d8341, 32'hc11e9ff8, 32'h427da796, 32'hc0a81cce, 32'h42754802, 32'h41a26306, 32'hc28f90e8};
test_label[1735] = '{32'hc11e9ff8};
test_output[1735] = '{32'h42d260d9};
/*############ DEBUG ############
test_input[13880:13887] = '{95.275099428, 70.7563567484, -9.91405463731, 63.4136587854, -5.25351633039, 61.3203205088, 20.2983507245, -71.7830194108};
test_label[1735] = '{-9.91405463731};
test_output[1735] = '{105.189154065};
############ END DEBUG ############*/
test_input[13888:13895] = '{32'hc299bdc9, 32'h41c4d197, 32'h427585b6, 32'hc186867b, 32'hc174ff50, 32'h4271411f, 32'h41557a12, 32'hc1c72205};
test_label[1736] = '{32'h4271411f};
test_output[1736] = '{32'h3fae6bce};
/*############ DEBUG ############
test_input[13888:13895] = '{-76.8706710296, 24.6023384877, 61.3805759081, -16.815663436, -15.3123324593, 60.3135952077, 13.3423027038, -24.8916118812};
test_label[1736] = '{60.3135952077};
test_output[1736] = '{1.36266496569};
############ END DEBUG ############*/
test_input[13896:13903] = '{32'h427863a1, 32'h42a1f6c4, 32'h41f44a2e, 32'h42c76000, 32'h428639ff, 32'h42a490d3, 32'hc1ea9041, 32'hc1453187};
test_label[1737] = '{32'h42a1f6c4};
test_output[1737] = '{32'h4195a4ef};
/*############ DEBUG ############
test_input[13896:13903] = '{62.0972920539, 80.9819637205, 30.5362196048, 99.6874982565, 67.1132746253, 82.2828594162, -29.3204361501, -12.3245914534};
test_label[1737] = '{80.9819637205};
test_output[1737] = '{18.7055345712};
############ END DEBUG ############*/
test_input[13904:13911] = '{32'hc2c34e72, 32'h421eb59e, 32'hc1ee7739, 32'hc28666b1, 32'hc2ba5c36, 32'hc13a62a7, 32'h429e84c2, 32'h42927467};
test_label[1738] = '{32'hc2ba5c36};
test_output[1738] = '{32'h432c7119};
/*############ DEBUG ############
test_input[13904:13911] = '{-97.6532154815, 39.6773594998, -29.8082134257, -67.2005698347, -93.1801008373, -11.6490853002, 79.2592944354, 73.2273460744};
test_label[1738] = '{-93.1801008373};
test_output[1738] = '{172.441793207};
############ END DEBUG ############*/
test_input[13912:13919] = '{32'hc28b11c3, 32'h42262065, 32'hc1958fa0, 32'h40f62250, 32'hc2824eb3, 32'h42150a23, 32'h4121c102, 32'h42988f4b};
test_label[1739] = '{32'h42262065};
test_output[1739] = '{32'h420afe32};
/*############ DEBUG ############
test_input[13912:13919] = '{-69.5346919316, 41.53163634, -18.6951288606, 7.69168854942, -65.1537111141, 37.2598996639, 10.1096210539, 76.2798726293};
test_label[1739] = '{41.53163634};
test_output[1739] = '{34.7482362893};
############ END DEBUG ############*/
test_input[13920:13927] = '{32'h429e7bde, 32'hc12ab22f, 32'h426b8341, 32'h42c76976, 32'hc2873735, 32'h418b275d, 32'h42ae4044, 32'h422e3e4d};
test_label[1740] = '{32'h418b275d};
test_output[1740] = '{32'h42a49f9f};
/*############ DEBUG ############
test_input[13920:13927] = '{79.2419274005, -10.6685015016, 58.8781771196, 99.7059747135, -67.6078277937, 17.3942195738, 87.1255190457, 43.5608388441};
test_label[1740] = '{17.3942195738};
test_output[1740] = '{82.3117585796};
############ END DEBUG ############*/
test_input[13928:13935] = '{32'h42aeb59d, 32'hc120a3c0, 32'hc2ba1fc8, 32'h423224e3, 32'hc2a5ed75, 32'h424d2657, 32'h42acd5ba, 32'h406d5f96};
test_label[1741] = '{32'h424d2657};
test_output[1741] = '{32'h42119758};
/*############ DEBUG ############
test_input[13928:13935] = '{87.3547150535, -10.0399781196, -93.062072, 44.5360215595, -82.9637859833, 51.2874408853, 86.4174375657, 3.70895908246};
test_label[1741] = '{51.2874408853};
test_output[1741] = '{36.397794997};
############ END DEBUG ############*/
test_input[13936:13943] = '{32'h42262b4e, 32'hc2a61fa1, 32'h4188b741, 32'h42a7c85d, 32'h42b99349, 32'h427a0daa, 32'hc2b5a52c, 32'h4288b7c6};
test_label[1742] = '{32'h42262b4e};
test_output[1742] = '{32'h424cfb69};
/*############ DEBUG ############
test_input[13936:13943] = '{41.5422884738, -83.0617720893, 17.0894788729, 83.8913309388, 92.7876680502, 62.5133456501, -90.8225982162, 68.3589317587};
test_label[1742] = '{41.5422884738};
test_output[1742] = '{51.2455164564};
############ END DEBUG ############*/
test_input[13944:13951] = '{32'hc2a0136e, 32'hc2c20b4c, 32'h428a45d2, 32'h42957f3d, 32'hc289be5f, 32'hc1a8476a, 32'hc29dfa5b, 32'hc26feb39};
test_label[1743] = '{32'h42957f3d};
test_output[1743] = '{32'h3b6efb4f};
/*############ DEBUG ############
test_input[13944:13951] = '{-80.0379515772, -97.0220647775, 69.1363672748, 74.7485114795, -68.8718182226, -21.034870269, -78.9889743837, -59.9797109066};
test_label[1743] = '{74.7485114795};
test_output[1743] = '{0.00364657085699};
############ END DEBUG ############*/
test_input[13952:13959] = '{32'h424b0f91, 32'h42af4fc8, 32'h422e77d8, 32'hc2a4a95d, 32'h41c390a1, 32'hc2c390c2, 32'h4229f99e, 32'h4295f8ac};
test_label[1744] = '{32'hc2a4a95d};
test_output[1744] = '{32'h4329fc93};
/*############ DEBUG ############
test_input[13952:13959] = '{50.7652034292, 87.6558260455, 43.6170354572, -82.3307865103, 24.4456201243, -97.7827322391, 42.4937658856, 74.985686539};
test_label[1744] = '{-82.3307865103};
test_output[1744] = '{169.986615699};
############ END DEBUG ############*/
test_input[13960:13967] = '{32'hc2540a7c, 32'hc24098a7, 32'h424383c3, 32'hc228a4bc, 32'hc1b27e65, 32'h425c8252, 32'hc1e1a3a6, 32'h421fee5e};
test_label[1745] = '{32'h425c8252};
test_output[1745] = '{32'h3afd2cf5};
/*############ DEBUG ############
test_input[13960:13967] = '{-53.0102389098, -48.1490741135, 48.878674472, -42.1608748426, -22.3117169163, 55.1272641681, -28.2049065242, 39.9827807864};
test_label[1745] = '{55.1272641681};
test_output[1745] = '{0.00193157663707};
############ END DEBUG ############*/
test_input[13968:13975] = '{32'hc0f1cbdb, 32'hc2c4a3ba, 32'h42014d99, 32'h42800043, 32'h428c3f1e, 32'h4286bce5, 32'h41d9647b, 32'h4258cc53};
test_label[1746] = '{32'h4258cc53};
test_output[1746] = '{32'h417fccd9};
/*############ DEBUG ############
test_input[13968:13975] = '{-7.55613490258, -98.3197776376, 32.3257771061, 64.0005129247, 70.1232788928, 67.3689357632, 27.1740636078, 54.1995335022};
test_label[1746] = '{54.1995335022};
test_output[1746] = '{15.9875117274};
############ END DEBUG ############*/
test_input[13976:13983] = '{32'h421efa4d, 32'hc22354b1, 32'hc2c1e13c, 32'hbfe6af4f, 32'h4286a609, 32'h41fd76bd, 32'hc2b6f56f, 32'h42c0610b};
test_label[1747] = '{32'h4286a609};
test_output[1747] = '{32'h41e6ec09};
/*############ DEBUG ############
test_input[13976:13983] = '{39.7444338849, -40.8327051513, -96.9399100755, -1.80222505123, 67.3242852831, 31.682978229, -91.4793653059, 96.1895363405};
test_label[1747] = '{67.3242852831};
test_output[1747] = '{28.8652510574};
############ END DEBUG ############*/
test_input[13984:13991] = '{32'h41ba8f80, 32'hc1372fe9, 32'h42b0cdb2, 32'hc299a8ac, 32'hc154a81d, 32'h429ebcaf, 32'h42a514c4, 32'h425bb277};
test_label[1748] = '{32'h425bb277};
test_output[1748] = '{32'h4205ebf4};
/*############ DEBUG ############
test_input[13984:13991] = '{23.3200692332, -11.4491971572, 88.4017450339, -76.8294364718, -13.2910431246, 79.3685224543, 82.5405597357, 54.9242833294};
test_label[1748] = '{54.9242833294};
test_output[1748] = '{33.4804245541};
############ END DEBUG ############*/
test_input[13992:13999] = '{32'h42127a0f, 32'h42429b08, 32'h42c6a25d, 32'hc272ff27, 32'h42346a24, 32'h41b2f458, 32'hc123c76d, 32'h42024c3c};
test_label[1749] = '{32'h41b2f458};
test_output[1749] = '{32'h4299e546};
/*############ DEBUG ############
test_input[13992:13999] = '{36.6191975962, 48.6513994764, 99.3171122454, -60.7491716319, 45.10365382, 22.3693088671, -10.2361875348, 32.5744485042};
test_label[1749] = '{22.3693088671};
test_output[1749] = '{76.9478033784};
############ END DEBUG ############*/
test_input[14000:14007] = '{32'h428194d5, 32'hc29ec52e, 32'hbf43b4cb, 32'h429d2b85, 32'hc2b199cc, 32'hc2681636, 32'h427bc921, 32'hc1bc91fb};
test_label[1750] = '{32'hc1bc91fb};
test_output[1750] = '{32'h42cc5004};
/*############ DEBUG ############
test_input[14000:14007] = '{64.7906899967, -79.3851154299, -0.764477425704, 78.5849999685, -88.8003854379, -58.0216896218, 62.9464167188, -23.5712786035};
test_label[1750] = '{-23.5712786035};
test_output[1750] = '{102.156279755};
############ END DEBUG ############*/
test_input[14008:14015] = '{32'hc1c6567e, 32'h41c70f74, 32'hc09c2cdb, 32'h42bd417a, 32'hc1bc30f2, 32'h4214c255, 32'hc2a56d95, 32'hc2aa59a8};
test_label[1751] = '{32'hc1c6567e};
test_output[1751] = '{32'h42eed71a};
/*############ DEBUG ############
test_input[14008:14015] = '{-24.7922315826, 24.8825460201, -4.8804756023, 94.6278852939, -23.5238987193, 37.189778506, -82.7140251117, -85.1751080185};
test_label[1751] = '{-24.7922315826};
test_output[1751] = '{119.420116877};
############ END DEBUG ############*/
test_input[14016:14023] = '{32'h42a53ef1, 32'h42aefca3, 32'hc1b2326e, 32'hc1fef9c9, 32'h425357e9, 32'hc2be9263, 32'h4259f904, 32'h423c1ee1};
test_label[1752] = '{32'hc1fef9c9};
test_output[1752] = '{32'h42eebeff};
/*############ DEBUG ############
test_input[14016:14023] = '{82.6229348578, 87.4934307869, -22.2746232664, -31.8719658928, 52.8358489592, -95.2859104112, 54.4931805702, 47.0301567113};
test_label[1752] = '{-31.8719658928};
test_output[1752] = '{119.373036979};
############ END DEBUG ############*/
test_input[14024:14031] = '{32'hc29abf70, 32'h428dd29c, 32'hc1ec2928, 32'hc23e8cb1, 32'hc2aba517, 32'hc2be707f, 32'hc218267b, 32'hc26dc140};
test_label[1753] = '{32'hc2be707f};
test_output[1753] = '{32'h4326218e};
/*############ DEBUG ############
test_input[14024:14031] = '{-77.3738993783, 70.911348367, -29.5200960403, -47.6373948604, -85.8224426074, -95.2197218957, -38.0375768313, -59.438721696};
test_label[1753] = '{-95.2197218957};
test_output[1753] = '{166.131070263};
############ END DEBUG ############*/
test_input[14032:14039] = '{32'h4285566d, 32'h42a5dabb, 32'h41a99df5, 32'hc284ca4f, 32'hc1e5e5e3, 32'hc15057bc, 32'h42a0a1ad, 32'hc2695031};
test_label[1754] = '{32'hc284ca4f};
test_output[1754] = '{32'h431564a9};
/*############ DEBUG ############
test_input[14032:14039] = '{66.6687997074, 82.9272060739, 21.202127304, -66.39513228, -28.7372488055, -13.0214195783, 80.3157759626, -58.3283134611};
test_label[1754] = '{-66.39513228};
test_output[1754] = '{149.393197057};
############ END DEBUG ############*/
test_input[14040:14047] = '{32'h42af0584, 32'h4299578d, 32'hc27f7ef8, 32'hc26e764e, 32'h42115c80, 32'h40622ceb, 32'h40bb9a0d, 32'hc2987432};
test_label[1755] = '{32'hc26e764e};
test_output[1755] = '{32'h43132057};
/*############ DEBUG ############
test_input[14040:14047] = '{87.5107743071, 76.6709973008, -63.8739947804, -59.6155317031, 36.3403311962, 3.53399156645, 5.86255513015, -76.226940877};
test_label[1755] = '{-59.6155317031};
test_output[1755] = '{147.126325614};
############ END DEBUG ############*/
test_input[14048:14055] = '{32'h412e1c7c, 32'h42b6dac2, 32'hc1222880, 32'h425b8664, 32'hc282ee36, 32'h42c1ab60, 32'hc20da91b, 32'h42a203a6};
test_label[1756] = '{32'hc1222880};
test_output[1756] = '{32'h42d5f2bb};
/*############ DEBUG ############
test_input[14048:14055] = '{10.8819540827, 91.4272632371, -10.1348881182, 54.8812404876, -65.4652537336, 96.8347200038, -35.4151417689, 81.0071230695};
test_label[1756] = '{-10.1348881182};
test_output[1756] = '{106.974081263};
############ END DEBUG ############*/
test_input[14056:14063] = '{32'h40327b19, 32'h4275a7f8, 32'hc284af3a, 32'h421e2a59, 32'hc140977d, 32'hc2a744dc, 32'hc239be7d, 32'h408db701};
test_label[1757] = '{32'h408db701};
test_output[1757] = '{32'h4263f118};
/*############ DEBUG ############
test_input[14056:14063] = '{2.78876321337, 61.4140325288, -66.3422367227, 39.5413540861, -12.0369842835, -83.6344875688, -46.4360236609, 4.42858917268};
test_label[1757] = '{4.42858917268};
test_output[1757] = '{56.9854433565};
############ END DEBUG ############*/
test_input[14064:14071] = '{32'hc282dac2, 32'hc2c42a67, 32'h4231eaa8, 32'h42a400a3, 32'hc24c1ddf, 32'h41502900, 32'hc28d9340, 32'h40831fb4};
test_label[1758] = '{32'hc24c1ddf};
test_output[1758] = '{32'h430507c9};
/*############ DEBUG ############
test_input[14064:14071] = '{-65.4272577324, -98.0828139647, 44.479156067, 82.0012443768, -51.0291718244, 13.0100099932, -70.787595494, 4.09762024447};
test_label[1758] = '{-51.0291718244};
test_output[1758] = '{133.030416201};
############ END DEBUG ############*/
test_input[14072:14079] = '{32'h42b3b7c8, 32'hc231c64f, 32'h42bfd1a1, 32'hc27578e1, 32'h41600cc2, 32'h428e9838, 32'hc1f1fb50, 32'h429ecacc};
test_label[1759] = '{32'hc1f1fb50};
test_output[1759] = '{32'h42fc51aa};
/*############ DEBUG ############
test_input[14072:14079] = '{89.8589504427, -44.4436613106, 95.9094324743, -61.3680476453, 14.0031151543, 71.2972998928, -30.2477115353, 79.3960849545};
test_label[1759] = '{-30.2477115353};
test_output[1759] = '{126.15949803};
############ END DEBUG ############*/
test_input[14080:14087] = '{32'hc2582a0a, 32'hc1992c63, 32'hc2ba4488, 32'h427f9446, 32'hc25b06cf, 32'hc2972a82, 32'hc26313a1, 32'h41eb27d0};
test_label[1760] = '{32'hc2582a0a};
test_output[1760] = '{32'h42ebdf28};
/*############ DEBUG ############
test_input[14080:14087] = '{-54.0410527514, -19.1466728917, -93.1338483789, 63.8947979844, -54.7566478264, -75.5830254495, -56.7691670214, 29.3944390325};
test_label[1760] = '{-54.0410527514};
test_output[1760] = '{117.935850736};
############ END DEBUG ############*/
test_input[14088:14095] = '{32'hc0362ef2, 32'hc2891217, 32'h42b965c0, 32'hc24a28fc, 32'h42332035, 32'h42972df8, 32'h42269225, 32'hc2964fa9};
test_label[1761] = '{32'h42332035};
test_output[1761] = '{32'h423fab4b};
/*############ DEBUG ############
test_input[14088:14095] = '{-2.84661522069, -68.5353349049, 92.6987311545, -50.5400245136, 44.7814520048, 75.5897842559, 41.6427183118, -75.1555871698};
test_label[1761] = '{44.7814520048};
test_output[1761] = '{47.9172791868};
############ END DEBUG ############*/
test_input[14096:14103] = '{32'hc013775f, 32'h428b264f, 32'h429fb7a5, 32'h42743197, 32'hc2a2d453, 32'h42881759, 32'h4247028f, 32'hc285bc88};
test_label[1762] = '{32'h42881759};
test_output[1762] = '{32'h413d028b};
/*############ DEBUG ############
test_input[14096:14103] = '{-2.30416088964, 69.5748179216, 79.8586790264, 61.0484258872, -81.4146964229, 68.0455996975, 49.7525002564, -66.8682241608};
test_label[1762] = '{68.0455996975};
test_output[1762] = '{11.8131209221};
############ END DEBUG ############*/
test_input[14104:14111] = '{32'hc0e40ba7, 32'h42c74eb6, 32'hc21eac34, 32'h4219db92, 32'h429fb052, 32'hc201b087, 32'hc2bada52, 32'h42bf3753};
test_label[1763] = '{32'hc2bada52};
test_output[1763] = '{32'h434118f5};
/*############ DEBUG ############
test_input[14104:14111] = '{-7.12642244954, 99.6537360549, -39.6681687296, 38.4644230642, 79.8443751377, -32.4223883988, -93.4264101151, 95.6080546774};
test_label[1763] = '{-93.4264101151};
test_output[1763] = '{193.097492627};
############ END DEBUG ############*/
test_input[14112:14119] = '{32'hc2047db8, 32'h411b1be1, 32'h42a98eab, 32'h42be2802, 32'hc22ffcf2, 32'hc2876968, 32'hc2adcfa9, 32'h41f581b2};
test_label[1764] = '{32'hc2047db8};
test_output[1764] = '{32'h43003371};
/*############ DEBUG ############
test_input[14112:14119] = '{-33.1227740641, 9.69430670774, 84.778648709, 95.07813821, -43.9970177491, -67.7058731794, -86.9055866328, 30.6883283777};
test_label[1764] = '{-33.1227740641};
test_output[1764] = '{128.200945924};
############ END DEBUG ############*/
test_input[14120:14127] = '{32'hc23deccd, 32'h40252f41, 32'hc288978d, 32'hc291d975, 32'hc210d90a, 32'hc0eaf0ed, 32'h41e1a1a7, 32'hc2ad8908};
test_label[1765] = '{32'hc288978d};
test_output[1765] = '{32'h42c0fff6};
/*############ DEBUG ############
test_input[14120:14127] = '{-47.4812491001, 2.58100906888, -68.2959948299, -72.9247205233, -36.2119508228, -7.34190987325, 28.2039316685, -86.7676400213};
test_label[1765] = '{-68.2959948299};
test_output[1765] = '{96.4999264984};
############ END DEBUG ############*/
test_input[14128:14135] = '{32'hc234c4c4, 32'h4294dcfe, 32'h429b0eeb, 32'h425fa97c, 32'h42905cc4, 32'h42968cdf, 32'hc28329fd, 32'hc2245f21};
test_label[1766] = '{32'h42905cc4};
test_output[1766] = '{32'h40afbe2d};
/*############ DEBUG ############
test_input[14128:14135] = '{-45.1921534269, 74.4316277436, 77.5291380398, 55.915511877, 72.1811850774, 75.2751385053, -65.5820057424, -41.092900798};
test_label[1766] = '{72.1811850774};
test_output[1766] = '{5.49196490501};
############ END DEBUG ############*/
test_input[14136:14143] = '{32'h422c6456, 32'hc2198cf0, 32'h422425c0, 32'h42612806, 32'hc20227e8, 32'h42a76b33, 32'hbe93bbcc, 32'h42afa363};
test_label[1767] = '{32'hc2198cf0};
test_output[1767] = '{32'h42fc7231};
/*############ DEBUG ############
test_input[14136:14143] = '{43.097985167, -38.3876343363, 41.0368649242, 56.2890853855, -32.5389692033, 83.7093760345, -0.288542146404, 87.8191154667};
test_label[1767] = '{-38.3876343363};
test_output[1767] = '{126.223028631};
############ END DEBUG ############*/
test_input[14144:14151] = '{32'h419c68cd, 32'h42a76108, 32'h42a9f9c9, 32'h40a52fc6, 32'h42412e8e, 32'h41d44085, 32'hc2303678, 32'h426e334a};
test_label[1768] = '{32'h42a9f9c9};
test_output[1768] = '{32'h3e77275d};
/*############ DEBUG ############
test_input[14144:14151] = '{19.5511731003, 83.6895107938, 84.9878652688, 5.16208192134, 48.295463416, 26.5315028654, -44.0531923118, 59.5500873649};
test_label[1768] = '{84.9878652688};
test_output[1768] = '{0.241361095661};
############ END DEBUG ############*/
test_input[14152:14159] = '{32'hc2163561, 32'hc210a704, 32'hc29a8aad, 32'hc1d65c78, 32'h42c33e58, 32'h4251ad2a, 32'hc2114685, 32'hc20ca22c};
test_label[1769] = '{32'h42c33e58};
test_output[1769] = '{32'h80000000};
/*############ DEBUG ############
test_input[14152:14159] = '{-37.5521280328, -36.1631000439, -77.2708478704, -26.7951508202, 97.6217643671, 52.4191045084, -36.3188665022, -35.1583726625};
test_label[1769] = '{97.6217643671};
test_output[1769] = '{-0.0};
############ END DEBUG ############*/
test_input[14160:14167] = '{32'hc23eb9e2, 32'h41953526, 32'h425118d9, 32'hc2902ad8, 32'h421996f5, 32'h42bdea1b, 32'h429f1d83, 32'hc1c7902a};
test_label[1770] = '{32'h42bdea1b};
test_output[1770] = '{32'h345c433b};
/*############ DEBUG ############
test_input[14160:14167] = '{-47.6815279163, 18.6509513111, 52.2742651269, -72.0836762632, 38.3974191515, 94.9572363329, 79.5576415964, -24.9453926745};
test_label[1770] = '{94.9572363329};
test_output[1770] = '{2.05135553601e-07};
############ END DEBUG ############*/
test_input[14168:14175] = '{32'hc26a2172, 32'hc295cb95, 32'h42beb94c, 32'h4263cd7b, 32'hc27e5cc7, 32'h41ffe7b7, 32'hc22f50a6, 32'hc23c6cc0};
test_label[1771] = '{32'hc23c6cc0};
test_output[1771] = '{32'h430e77d6};
/*############ DEBUG ############
test_input[14168:14175] = '{-58.5326628564, -74.8976185277, 95.3619051165, 56.9506660916, -63.5906035923, 31.9881423221, -43.8287590889, -47.1062012191};
test_label[1771] = '{-47.1062012191};
test_output[1771] = '{142.468106336};
############ END DEBUG ############*/
test_input[14176:14183] = '{32'h42b4b7e2, 32'h40f0abe7, 32'hc1ce5928, 32'hc1ec8b12, 32'h42c3f794, 32'hc2c4acf2, 32'h413e8a0f, 32'h4282811c};
test_label[1772] = '{32'hc2c4acf2};
test_output[1772] = '{32'h43445263};
/*############ DEBUG ############
test_input[14176:14183] = '{90.3591469383, 7.52098430874, -25.7935333215, -29.5679045586, 97.9835514409, -98.3377863748, 11.9087058223, 65.2521646182};
test_label[1772] = '{-98.3377863748};
test_output[1772] = '{196.321826082};
############ END DEBUG ############*/
test_input[14184:14191] = '{32'hc29892af, 32'h42713d81, 32'h413f025e, 32'h429d32ab, 32'hc297cb91, 32'h42a17e05, 32'hc27cbd01, 32'h4211a11f};
test_label[1773] = '{32'h4211a11f};
test_output[1773] = '{32'h4231cc0c};
/*############ DEBUG ############
test_input[14184:14191] = '{-76.2864876901, 60.3100605026, 11.9380780575, 78.5989582038, -75.8975901835, 80.7461315162, -63.1845723014, 36.4073458357};
test_label[1773] = '{36.4073458357};
test_output[1773] = '{44.4492655702};
############ END DEBUG ############*/
test_input[14192:14199] = '{32'h42984518, 32'hc278b625, 32'h4109667e, 32'hc0dcda5f, 32'hc23452b6, 32'h4264ddbc, 32'h41b420cf, 32'hc0c3e339};
test_label[1774] = '{32'hc0dcda5f};
test_output[1774] = '{32'h42a612be};
/*############ DEBUG ############
test_input[14192:14199] = '{76.134950551, -62.1778757926, 8.58752208349, -6.9016564093, -45.0807715336, 57.2165373667, 22.5160205433, -6.12148706517};
test_label[1774] = '{-6.9016564093};
test_output[1774] = '{83.0366069663};
############ END DEBUG ############*/
test_input[14200:14207] = '{32'h42b63989, 32'h41874f30, 32'hc17f92b5, 32'h4249520e, 32'hc22f896d, 32'h4264119b, 32'hc264585e, 32'hc2b45f88};
test_label[1775] = '{32'hc22f896d};
test_output[1775] = '{32'h4306ff20};
/*############ DEBUG ############
test_input[14200:14207] = '{91.1123717273, 16.9136655732, -15.9733173328, 50.3301298939, -43.8842032412, 57.0171929545, -57.0862962104, -90.1865859594};
test_label[1775] = '{-43.8842032412};
test_output[1775] = '{134.996574968};
############ END DEBUG ############*/
test_input[14208:14215] = '{32'hc136a4dd, 32'hc04c29c6, 32'h422dc3ea, 32'h42af52f8, 32'h4241508a, 32'hc2c0d8c2, 32'h42ad2d15, 32'h423036c5};
test_label[1776] = '{32'h42ad2d15};
test_output[1776] = '{32'h3faf1708};
/*############ DEBUG ############
test_input[14208:14215] = '{-11.4152501584, -3.19004953385, 43.4413239854, 87.6620451323, 48.3286506147, -96.4233579845, 86.5880474946, 44.0534854232};
test_label[1776] = '{86.5880474946};
test_output[1776] = '{1.36789040691};
############ END DEBUG ############*/
test_input[14216:14223] = '{32'h429b4592, 32'h42853bf0, 32'h41911200, 32'h410b7b39, 32'hc110c8bb, 32'h42b1fde6, 32'hc2b81f11, 32'h42079729};
test_label[1777] = '{32'h42853bf0};
test_output[1777] = '{32'h41b307db};
/*############ DEBUG ############
test_input[14216:14223] = '{77.6358772616, 66.6170684347, 18.1337896336, 8.71758321342, -9.04900681491, 88.9958926102, -92.0606782642, 33.8976184974};
test_label[1777] = '{66.6170684347};
test_output[1777] = '{22.3788358279};
############ END DEBUG ############*/
test_input[14224:14231] = '{32'hc2167075, 32'hc2c2067a, 32'hc13f35d8, 32'h41a4c382, 32'h3febc870, 32'h42ab8736, 32'h41940b07, 32'hc2c6194b};
test_label[1778] = '{32'h41940b07};
test_output[1778] = '{32'h42868474};
/*############ DEBUG ############
test_input[14224:14231] = '{-37.60982182, -97.0126461031, -11.9506451253, 20.5954637227, 1.84205437912, 85.7640836361, 18.505384416, -99.0493977535};
test_label[1778] = '{18.505384416};
test_output[1778] = '{67.2586992202};
############ END DEBUG ############*/
test_input[14232:14239] = '{32'hc28de06e, 32'h42b6cb76, 32'hc2b239e9, 32'h42bcc39d, 32'hc1b6bf5c, 32'hc295cda9, 32'hc254127b, 32'h4116ca72};
test_label[1779] = '{32'hc28de06e};
test_output[1779] = '{32'h43255ea6};
/*############ DEBUG ############
test_input[14232:14239] = '{-70.9383425846, 91.3973871055, -89.1131058351, 94.3820579848, -22.8434372421, -74.901678368, -53.018047847, 9.4244249003};
test_label[1779] = '{-70.9383425846};
test_output[1779] = '{165.36972025};
############ END DEBUG ############*/
test_input[14240:14247] = '{32'h4247ec87, 32'hc2835595, 32'h425e44e1, 32'hc22c0937, 32'h3fa04884, 32'h409f35f7, 32'h42835a40, 32'h42095100};
test_label[1780] = '{32'h409f35f7};
test_output[1780] = '{32'h4272cdcd};
/*############ DEBUG ############
test_input[14240:14247] = '{49.9809852997, -65.6671533775, 55.5672657452, -43.0089981216, 1.25221303853, 4.97533742466, 65.6762726496, 34.3291022511};
test_label[1780] = '{4.97533742466};
test_output[1780] = '{60.700976088};
############ END DEBUG ############*/
test_input[14248:14255] = '{32'h428a4362, 32'hc2c41ae8, 32'h3f1528f8, 32'hc2060fb3, 32'h419cf401, 32'hc2bb9cd2, 32'h41703079, 32'hc0fe9c19};
test_label[1781] = '{32'h428a4362};
test_output[1781] = '{32'h80000000};
/*############ DEBUG ############
test_input[14248:14255] = '{69.1316073434, -98.0525530602, 0.582656370214, -33.5153313007, 19.6191419448, -93.806286097, 15.0118340293, -7.95655468705};
test_label[1781] = '{69.1316073434};
test_output[1781] = '{-0.0};
############ END DEBUG ############*/
test_input[14256:14263] = '{32'h42c42d9d, 32'h4239cf9e, 32'hc236349c, 32'h41b52671, 32'h4122ef96, 32'hc1c238af, 32'hc2688cda, 32'h421cde72};
test_label[1782] = '{32'h4239cf9e};
test_output[1782] = '{32'h424e8b9c};
/*############ DEBUG ############
test_input[14256:14263] = '{98.0890887407, 46.452750194, -45.5513773004, 22.6437706349, 10.1834929184, -24.2776781186, -58.1375495635, 39.2172322004};
test_label[1782] = '{46.452750194};
test_output[1782] = '{51.6363385467};
############ END DEBUG ############*/
test_input[14264:14271] = '{32'hc09dab48, 32'h424d30d4, 32'h4274162f, 32'hc10f44bc, 32'hc21bb3c0, 32'h421df442, 32'h411ed306, 32'h42b335fd};
test_label[1783] = '{32'h4274162f};
test_output[1783] = '{32'h41e4ab96};
/*############ DEBUG ############
test_input[14264:14271] = '{-4.92715838305, 51.2976841213, 61.0216635498, -8.95428047821, -38.9255370681, 39.4885347254, 9.92651943511, 89.6054456685};
test_label[1783] = '{61.0216635498};
test_output[1783] = '{28.5837821187};
############ END DEBUG ############*/
test_input[14272:14279] = '{32'hc2a88c81, 32'h4140d0d6, 32'hc25e44e3, 32'h41db9569, 32'hc275fac3, 32'hc2c3585e, 32'h4266305e, 32'h402c3447};
test_label[1784] = '{32'hc2a88c81};
test_output[1784] = '{32'h430dd258};
/*############ DEBUG ############
test_input[14272:14279] = '{-84.2744224914, 12.0509854818, -55.5672729437, 27.447954421, -61.4948830289, -97.672589234, 57.547233313, 2.69069066376};
test_label[1784] = '{-84.2744224914};
test_output[1784] = '{141.821655804};
############ END DEBUG ############*/
test_input[14280:14287] = '{32'hc252d182, 32'hc2a1d63b, 32'hc2b77146, 32'hc1af3fb6, 32'h42945b5e, 32'h42b8991f, 32'hc0939c93, 32'hc1e7dd90};
test_label[1785] = '{32'h42b8991f};
test_output[1785] = '{32'h3267eb34};
/*############ DEBUG ############
test_input[14280:14287] = '{-52.7045962922, -80.9184213106, -91.7212348902, -21.9061088823, 74.1784484726, 92.2990654496, -4.61286300319, -28.9831845316};
test_label[1785] = '{92.2990654496};
test_output[1785] = '{1.34994487611e-08};
############ END DEBUG ############*/
test_input[14288:14295] = '{32'h419395d7, 32'hc2321cdf, 32'h428fb293, 32'h42bedf70, 32'hc1ba06c2, 32'h41b849e6, 32'h424d443c, 32'h418811b3};
test_label[1786] = '{32'hc2321cdf};
test_output[1786] = '{32'h430bf6f0};
/*############ DEBUG ############
test_input[14288:14295] = '{18.4481631449, -44.5281945283, 71.8487790901, 95.4364049992, -23.25330006, 23.0360827125, 51.3166345921, 17.0086423659};
test_label[1786] = '{-44.5281945283};
test_output[1786] = '{139.964599528};
############ END DEBUG ############*/
test_input[14296:14303] = '{32'hc142c85f, 32'h4130fa83, 32'hc2a1fd3f, 32'h41fd143c, 32'hc28866c7, 32'h4282f702, 32'h41184ac0, 32'hc2b80f63};
test_label[1787] = '{32'hc142c85f};
test_output[1787] = '{32'h429b500e};
/*############ DEBUG ############
test_input[14296:14303] = '{-12.1739182494, 11.0611603055, -80.9946221095, 31.6348803561, -68.2007387723, 65.4824349743, 9.51824966572, -92.0300515194};
test_label[1787] = '{-12.1739182494};
test_output[1787] = '{77.6563532237};
############ END DEBUG ############*/
test_input[14304:14311] = '{32'hc23d8790, 32'h42685b45, 32'hc275f5cc, 32'hc278f60d, 32'hc21cbdea, 32'h429e8fad, 32'hc29328a1, 32'hc08a4d14};
test_label[1788] = '{32'hc23d8790};
test_output[1788] = '{32'h42fd5375};
/*############ DEBUG ############
test_input[14304:14311] = '{-47.3823862901, 58.0891299336, -61.4900348279, -62.2402843213, -39.1854612631, 79.2806156881, -73.579356875, -4.32190910521};
test_label[1788] = '{-47.3823862901};
test_output[1788] = '{126.663001979};
############ END DEBUG ############*/
test_input[14312:14319] = '{32'hc16f0418, 32'hc2b62ad1, 32'hc1d086c8, 32'hc299721e, 32'hc2294f79, 32'hc2b00787, 32'hc25e97e1, 32'h40704664};
test_label[1789] = '{32'hc299721e};
test_output[1789] = '{32'h42a0f452};
/*############ DEBUG ############
test_input[14312:14319] = '{-14.9384992646, -91.0836227859, -26.0658106456, -76.7228887708, -42.3276092258, -88.0147008974, -55.6483181922, 3.75429635608};
test_label[1789] = '{-76.7228887708};
test_output[1789] = '{80.4771851345};
############ END DEBUG ############*/
test_input[14320:14327] = '{32'h418c0a17, 32'hc2a547b5, 32'hc27ca903, 32'h42908faa, 32'h42092f9e, 32'hc2c3c9bb, 32'hc20ed9b9, 32'hc28fae7d};
test_label[1790] = '{32'hc2a547b5};
test_output[1790] = '{32'h431aebb0};
/*############ DEBUG ############
test_input[14320:14327] = '{17.5049262995, -82.6400552105, -63.1650513432, 72.2805919296, 34.2964998517, -97.8940031155, -35.712619482, -71.8407957107};
test_label[1790] = '{-82.6400552105};
test_output[1790] = '{154.92064714};
############ END DEBUG ############*/
test_input[14328:14335] = '{32'h41c1465b, 32'h427b2762, 32'h41b13745, 32'h42653639, 32'hc22ba460, 32'h426df1b0, 32'hc2c26a1d, 32'hc26bb2cb};
test_label[1791] = '{32'h427b2762};
test_output[1791] = '{32'h3d245906};
/*############ DEBUG ############
test_input[14328:14335] = '{24.1593524481, 62.7884596324, 22.1519867546, 57.3029526891, -42.910521481, 59.486022011, -97.2072556311, -58.9246028286};
test_label[1791] = '{62.7884596324};
test_output[1791] = '{0.0401239610966};
############ END DEBUG ############*/
test_input[14336:14343] = '{32'h41e1c350, 32'hc26df2b8, 32'hc1f3664a, 32'hc2197432, 32'hc14f2906, 32'hc28fc1cc, 32'hc2c6d026, 32'h421aa649};
test_label[1792] = '{32'hc26df2b8};
test_output[1792] = '{32'h42c44c84};
/*############ DEBUG ############
test_input[14336:14343] = '{28.2203674954, -59.4870307075, -30.4249461925, -38.3634723529, -12.9475154356, -71.8785074731, -99.4065415466, 38.662387808};
test_label[1792] = '{-59.4870307075};
test_output[1792] = '{98.1494476953};
############ END DEBUG ############*/
test_input[14344:14351] = '{32'hc2c5a8da, 32'h42b6bc9d, 32'hc2b149fd, 32'hc29ead4d, 32'h42ba838c, 32'h4202cb8d, 32'h429c1dc1, 32'hc29bf095};
test_label[1793] = '{32'hc2c5a8da};
test_output[1793] = '{32'h43403a44};
/*############ DEBUG ############
test_input[14344:14351] = '{-98.8297869822, 91.3683822387, -88.6445088627, -79.3384760224, 93.2569254382, 32.6987799705, 78.0581162777, -77.9698884209};
test_label[1793] = '{-98.8297869822};
test_output[1793] = '{192.227597472};
############ END DEBUG ############*/
test_input[14352:14359] = '{32'hc16fa303, 32'hc1b8d729, 32'h42894fc6, 32'h4225e928, 32'h427290e2, 32'hc2976c09, 32'hc2a47ed0, 32'h42a57f1f};
test_label[1794] = '{32'hc1b8d729};
test_output[1794] = '{32'h42d3b4e9};
/*############ DEBUG ############
test_input[14352:14359] = '{-14.9772982359, -23.1050587862, 68.6558065682, 41.4776930231, 60.6414867841, -75.7110072339, -82.2476826105, 82.7482829408};
test_label[1794] = '{-23.1050587862};
test_output[1794] = '{105.853342485};
############ END DEBUG ############*/
test_input[14360:14367] = '{32'h4271e575, 32'hc191dddd, 32'hc295e2e7, 32'hc2bcd09a, 32'hbfabed8a, 32'hc2970524, 32'hc26fa71c, 32'h42366008};
test_label[1795] = '{32'hbfabed8a};
test_output[1795] = '{32'h427744e2};
/*############ DEBUG ############
test_input[14360:14367] = '{60.4740797392, -18.2333324174, -74.9431650376, -94.4074248521, -1.34318660417, -75.5100429082, -59.9131912274, 45.593781154};
test_label[1795] = '{-1.34318660417};
test_output[1795] = '{61.8172666881};
############ END DEBUG ############*/
test_input[14368:14375] = '{32'hc2328c7d, 32'hc2527098, 32'h40bf027c, 32'hc2a52a65, 32'h428ea541, 32'hc21ce9a1, 32'hc2084c3a, 32'h428995c8};
test_label[1796] = '{32'hc2328c7d};
test_output[1796] = '{32'h42e812bb};
/*############ DEBUG ############
test_input[14368:14375] = '{-44.6371939085, -52.6099556911, 5.96905315679, -82.5827996455, 71.3227614069, -39.2281547561, -34.0744385058, 68.7925430082};
test_label[1796] = '{-44.6371939085};
test_output[1796] = '{116.036584472};
############ END DEBUG ############*/
test_input[14376:14383] = '{32'h420abfa0, 32'h42075ceb, 32'hc1ea8e6d, 32'hc1d0fbf7, 32'h42a95376, 32'hc24d7919, 32'hc12db400, 32'hc2b7ff74};
test_label[1797] = '{32'hc1d0fbf7};
test_output[1797] = '{32'h42dd9274};
/*############ DEBUG ############
test_input[14376:14383] = '{34.687132774, 33.8407385322, -29.3195439128, -26.1230288235, 84.6630119636, -51.3682611915, -10.8564456631, -91.9989336919};
test_label[1797] = '{-26.1230288235};
test_output[1797] = '{110.786040787};
############ END DEBUG ############*/
test_input[14384:14391] = '{32'h42b4b0e8, 32'h41fc93b3, 32'h41b831b0, 32'h424ec3f0, 32'hc2b48e57, 32'h4210bea3, 32'hc1caa5b7, 32'hc281038c};
test_label[1798] = '{32'h4210bea3};
test_output[1798] = '{32'h4258a32e};
/*############ DEBUG ############
test_input[14384:14391] = '{90.3455211511, 31.5721183669, 23.0242620078, 51.6913467175, -90.2780100841, 36.186167765, -25.3309160817, -64.5069258283};
test_label[1798] = '{36.186167765};
test_output[1798] = '{54.1593533861};
############ END DEBUG ############*/
test_input[14392:14399] = '{32'hc1c03592, 32'h42982e3d, 32'h429282ee, 32'h4291cb4e, 32'h42b1cc9d, 32'hc298461a, 32'h3fd4f102, 32'h42a725c3};
test_label[1799] = '{32'h3fd4f102};
test_output[1799] = '{32'h42ae7b56};
/*############ DEBUG ############
test_input[14392:14399] = '{-24.0261568247, 76.0903126718, 73.2557217373, 72.8970800667, 88.8996371796, -76.1369156822, 1.6636049392, 83.5737527506};
test_label[1799] = '{1.6636049392};
test_output[1799] = '{87.2408874899};
############ END DEBUG ############*/
test_input[14400:14407] = '{32'h40611ecf, 32'hc29f9c54, 32'hc1626aff, 32'h422ed3e0, 32'h4223185a, 32'hc090a5fe, 32'h421284bc, 32'hc08698fa};
test_label[1800] = '{32'h40611ecf};
test_output[1800] = '{32'h4220f7e0};
/*############ DEBUG ############
test_input[14400:14407] = '{3.51750536414, -79.8053274379, -14.1511218623, 43.7069088735, 40.7737804313, -4.52026252415, 36.629623084, -4.20617370083};
test_label[1800] = '{3.51750536414};
test_output[1800] = '{40.2420664605};
############ END DEBUG ############*/
test_input[14408:14415] = '{32'hc2be205f, 32'h42261288, 32'h41546fcf, 32'hc2087bd5, 32'hc2064bc2, 32'hc180545b, 32'h428a88e3, 32'hc1d5ebba};
test_label[1801] = '{32'h41546fcf};
test_output[1801] = '{32'h425ff5d1};
/*############ DEBUG ############
test_input[14408:14415] = '{-95.0632217165, 41.5180969301, 13.2772969307, -34.1209309655, -33.5739840002, -16.0411887661, 69.2673536444, -26.7401009692};
test_label[1801] = '{13.2772969307};
test_output[1801] = '{55.9900567137};
############ END DEBUG ############*/
test_input[14416:14423] = '{32'h420a8fa4, 32'hc23efe1e, 32'hc28c6cba, 32'hc283daa1, 32'hc21381a3, 32'hc2571b55, 32'h428eb62a, 32'hc115f5cb};
test_label[1802] = '{32'h428eb62a};
test_output[1802] = '{32'h25000000};
/*############ DEBUG ############
test_input[14416:14423] = '{34.6402733962, -47.7481599573, -70.2123589174, -65.9270091296, -36.8765990829, -53.7766902858, 71.3557897287, -9.37250808431};
test_label[1802] = '{71.3557897287};
test_output[1802] = '{1.11022302463e-16};
############ END DEBUG ############*/
test_input[14424:14431] = '{32'h4249dc16, 32'h4238263d, 32'h421f4686, 32'hc26dfc35, 32'hc246acab, 32'h42a45473, 32'h41028712, 32'h42a196d6};
test_label[1803] = '{32'hc246acab};
test_output[1803] = '{32'h43040f57};
/*############ DEBUG ############
test_input[14424:14431] = '{50.4649273899, 46.0373421523, 39.8188723414, -59.4962941612, -49.6686210961, 82.1649428871, 8.15797644812, 80.7945986365};
test_label[1803] = '{-49.6686210961};
test_output[1803] = '{132.059917974};
############ END DEBUG ############*/
test_input[14432:14439] = '{32'hc02bf3b8, 32'h42ace2fc, 32'hc21c5747, 32'h418d5498, 32'hc1ce0a16, 32'h425d3252, 32'hc2c38161, 32'h4255d81a};
test_label[1804] = '{32'h418d5498};
test_output[1804] = '{32'h42898dd6};
/*############ DEBUG ############
test_input[14432:14439] = '{-2.68675040479, 86.4433282151, -39.0852302454, 17.666305379, -25.7549243917, 55.2991404604, -97.7526935848, 53.4610375594};
test_label[1804] = '{17.666305379};
test_output[1804] = '{68.7770228361};
############ END DEBUG ############*/
test_input[14440:14447] = '{32'h425bfe7b, 32'hc18979cb, 32'h4021cc3c, 32'hc2be8314, 32'h42c1d77b, 32'hc29efcb5, 32'h428541f3, 32'h4216fc5f};
test_label[1805] = '{32'h428541f3};
test_output[1805] = '{32'h41f25622};
/*############ DEBUG ############
test_input[14440:14447] = '{54.9985171653, -17.1844687325, 2.52809038458, -95.2560118676, 96.9208624167, -79.4935721381, 66.6288047303, 37.7464571351};
test_label[1805] = '{66.6288047303};
test_output[1805] = '{30.2920576864};
############ END DEBUG ############*/
test_input[14448:14455] = '{32'hc0312e55, 32'h415c7416, 32'hc1f331f9, 32'hc2b27400, 32'h4225ff43, 32'hc2ba041e, 32'h4213be15, 32'h42b23e2c};
test_label[1806] = '{32'hc1f331f9};
test_output[1806] = '{32'h42ef0aaa};
/*############ DEBUG ############
test_input[14448:14455] = '{-2.76845290868, 13.778341748, -30.3994005232, -89.2265640393, 41.4992771256, -93.0080428539, 36.9356279081, 89.1214285356};
test_label[1806] = '{-30.3994005232};
test_output[1806] = '{119.520829059};
############ END DEBUG ############*/
test_input[14456:14463] = '{32'h42860fb3, 32'hc2a44235, 32'h42a456e9, 32'hc29e1de5, 32'h42091ed2, 32'hc28910f5, 32'hc2025229, 32'hc2016a2b};
test_label[1807] = '{32'hc2025229};
test_output[1807] = '{32'h42e57ffe};
/*############ DEBUG ############
test_input[14456:14463] = '{67.0306625866, -82.1293134991, 82.1697469125, -79.0583904562, 34.2800990883, -68.5331179079, -32.580234443, -32.3536812939};
test_label[1807] = '{-32.580234443};
test_output[1807] = '{114.749981622};
############ END DEBUG ############*/
test_input[14464:14471] = '{32'hc2946133, 32'hc211cdcd, 32'hc0d3b179, 32'hc2a954ce, 32'h42796692, 32'h4110d666, 32'h42adac88, 32'h41f0d724};
test_label[1808] = '{32'hc2946133};
test_output[1808] = '{32'h432106de};
/*############ DEBUG ############
test_input[14464:14471] = '{-74.1898456654, -36.4509779547, -6.61541424948, -84.6656353524, 62.3501679237, 9.05234304548, 86.836973549, 30.1050500553};
test_label[1808] = '{-74.1898456654};
test_output[1808] = '{161.026819214};
############ END DEBUG ############*/
test_input[14472:14479] = '{32'hc2485815, 32'hc1c7b403, 32'h41b7ab09, 32'hc2a82a33, 32'h41e6fad6, 32'h42c2a1bb, 32'hc247f86f, 32'h41c53e8d};
test_label[1809] = '{32'h41b7ab09};
test_output[1809] = '{32'h4294b6f9};
/*############ DEBUG ############
test_input[14472:14479] = '{-50.0860185576, -24.96289559, 22.9585128462, -84.0824178285, 28.8724784357, 97.3158813707, -49.9926100991, 24.6555416657};
test_label[1809] = '{22.9585128462};
test_output[1809] = '{74.3573685245};
############ END DEBUG ############*/
test_input[14480:14487] = '{32'hc236b0d3, 32'hc2c72bab, 32'h41ca4ebb, 32'hc275ed08, 32'hc2aac3ae, 32'h429d5235, 32'h42906bb2, 32'h4185ea11};
test_label[1810] = '{32'h42906bb2};
test_output[1810] = '{32'h40ce751b};
/*############ DEBUG ############
test_input[14480:14487] = '{-45.6726804337, -99.5852906655, 25.2884419076, -61.4814774269, -85.3821891889, 78.6605597357, 72.210343382, 16.7392893258};
test_label[1810] = '{72.210343382};
test_output[1810] = '{6.45179528685};
############ END DEBUG ############*/
test_input[14488:14495] = '{32'h40ce76fb, 32'h41b77522, 32'h425b5feb, 32'hc165021f, 32'h428c3827, 32'h41eb47ab, 32'hc2385e8d, 32'h424d749f};
test_label[1811] = '{32'h425b5feb};
test_output[1811] = '{32'h41744191};
/*############ DEBUG ############
test_input[14488:14495] = '{6.45202402221, 22.9321932955, 54.8436689053, -14.3130175122, 70.1096760852, 29.4099934578, -46.0923359437, 51.3638870366};
test_label[1811] = '{54.8436689053};
test_output[1811] = '{15.2660074216};
############ END DEBUG ############*/
test_input[14496:14503] = '{32'h42bb90df, 32'h4274c6e4, 32'hc1f05aa7, 32'h427102c1, 32'h41546651, 32'h42a2edf2, 32'hc2349637, 32'hc2691751};
test_label[1812] = '{32'h42a2edf2};
test_output[1812] = '{32'h41451766};
/*############ DEBUG ############
test_input[14496:14503] = '{93.7829476733, 61.1942288188, -30.0442643275, 60.252688036, 13.2749799527, 81.464739878, -45.1466943311, -58.2727709212};
test_label[1812] = '{81.464739878};
test_output[1812] = '{12.3182122649};
############ END DEBUG ############*/
test_input[14504:14511] = '{32'hc2872378, 32'h4243f226, 32'hc2963b6e, 32'h4280d804, 32'h42344979, 32'hc28b6be1, 32'hc228a08e, 32'hc24a991f};
test_label[1813] = '{32'h42344979};
test_output[1813] = '{32'h419acd20};
/*############ DEBUG ############
test_input[14504:14511] = '{-67.5692739045, 48.9864746343, -75.1160724386, 64.4219090129, 45.0717500124, -69.7107014171, -42.1567932132, -50.6495311238};
test_label[1813] = '{45.0717500124};
test_output[1813] = '{19.3501592024};
############ END DEBUG ############*/
test_input[14512:14519] = '{32'h42bffff1, 32'h42906360, 32'h427a0492, 32'h40b4b4b1, 32'h420cdcd8, 32'hc27f1bcd, 32'hc22f97ad, 32'h4262ffbe};
test_label[1814] = '{32'h42906360};
test_output[1814] = '{32'h41be7245};
/*############ DEBUG ############
test_input[14512:14519] = '{95.9998850791, 72.1940891914, 62.5044647218, 5.64705711441, 35.2156692325, -63.7771490987, -43.8981195045, 56.7497500823};
test_label[1814] = '{72.1940891914};
test_output[1814] = '{23.8057958878};
############ END DEBUG ############*/
test_input[14520:14527] = '{32'h418d6be4, 32'h42c63ae9, 32'hc281ae02, 32'hc234548c, 32'h42a1aaec, 32'hc2a25bcc, 32'hc16e4283, 32'h417c1045};
test_label[1815] = '{32'h42a1aaec};
test_output[1815] = '{32'h41923ff7};
/*############ DEBUG ############
test_input[14520:14527] = '{17.6776806706, 99.1150625542, -64.839856081, -45.0825658145, 80.8338304154, -81.1792898911, -14.8912380823, 15.7539725086};
test_label[1815] = '{80.8338304154};
test_output[1815] = '{18.2812321503};
############ END DEBUG ############*/
test_input[14528:14535] = '{32'hc2651066, 32'h42861349, 32'h41847b6c, 32'hc24925b3, 32'hc292a476, 32'hc24fa3f8, 32'hc1e401e3, 32'hc2a1033d};
test_label[1816] = '{32'hc2651066};
test_output[1816] = '{32'h42f89b7c};
/*############ DEBUG ############
test_input[14528:14535] = '{-57.2660141421, 67.0376682094, 16.5602637389, -50.2868171271, -73.321211, -51.9101272277, -28.5009206003, -80.5063260528};
test_label[1816] = '{-57.2660141421};
test_output[1816] = '{124.303682352};
############ END DEBUG ############*/
test_input[14536:14543] = '{32'hc16ae73b, 32'h42935516, 32'h41ae0ecc, 32'h422d1241, 32'hc1cd1c11, 32'hc1ba4415, 32'h42b03a82, 32'h429072ba};
test_label[1817] = '{32'h41ae0ecc};
test_output[1817] = '{32'h4284b6cf};
/*############ DEBUG ############
test_input[14536:14543] = '{-14.6814524175, 73.666184391, 21.7572255326, 43.2678247842, -25.6387040992, -23.2832435285, 88.1142714799, 72.2240729275};
test_label[1817] = '{21.7572255326};
test_output[1817] = '{66.3570466042};
############ END DEBUG ############*/
test_input[14544:14551] = '{32'h4250d3b9, 32'h421c6026, 32'hc291073b, 32'h429e2c83, 32'hc2570bfe, 32'hc27886d8, 32'hc19eebb9, 32'h414e8ac0};
test_label[1818] = '{32'h414e8ac0};
test_output[1818] = '{32'h42845b2b};
/*############ DEBUG ############
test_input[14544:14551] = '{52.2067601829, 39.0938953931, -72.5141244845, 79.0869333941, -53.7617107869, -62.1316825401, -19.8650993263, 12.9088745043};
test_label[1818] = '{12.9088745043};
test_output[1818] = '{66.1780588898};
############ END DEBUG ############*/
test_input[14552:14559] = '{32'hc09762be, 32'h429e1476, 32'h428f1825, 32'h41294ae6, 32'h419f9f7a, 32'hc1423e3b, 32'hc1df97e8, 32'hc26a0f15};
test_label[1819] = '{32'h429e1476};
test_output[1819] = '{32'h3a11fe7c};
/*############ DEBUG ############
test_input[14552:14559] = '{-4.73080345797, 79.0399634731, 71.5471587907, 10.5807856429, 19.9528689421, -12.1401925172, -27.949172843, -58.5147281542};
test_label[1819] = '{79.0399634731};
test_output[1819] = '{0.00055692322901};
############ END DEBUG ############*/
test_input[14560:14567] = '{32'h41a28055, 32'h427e5f2d, 32'hc1468bb8, 32'hc18c6485, 32'hc297f4cc, 32'hc2a5f109, 32'h41e248c2, 32'h42bd2a68};
test_label[1820] = '{32'h41a28055};
test_output[1820] = '{32'h42948a53};
/*############ DEBUG ############
test_input[14560:14567] = '{20.3126615137, 63.5929434305, -12.4091109248, -17.5490809546, -75.9781197924, -82.9707747584, 28.2855258114, 94.5828273428};
test_label[1820] = '{20.3126615137};
test_output[1820] = '{74.2701658291};
############ END DEBUG ############*/
test_input[14568:14575] = '{32'hc2c01502, 32'h42bbcbf5, 32'h41f64f7d, 32'h423dcd25, 32'h4117b4df, 32'hc2797a13, 32'hbe9d6aa7, 32'h425b5218};
test_label[1821] = '{32'hbe9d6aa7};
test_output[1821] = '{32'h42bc6960};
/*############ DEBUG ############
test_input[14568:14575] = '{-96.0410297239, 93.8983551279, 30.788812734, 47.450337578, 9.48165753577, -62.3692113, -0.30745432725, 54.8301700561};
test_label[1821] = '{-0.30745432725};
test_output[1821] = '{94.2058094551};
############ END DEBUG ############*/
test_input[14576:14583] = '{32'h42b1b2b9, 32'h4236c3e7, 32'h4247eeb8, 32'hc20f9f71, 32'h42143040, 32'hc26a4db3, 32'hc2c269e5, 32'h4287d34f};
test_label[1822] = '{32'h42b1b2b9};
test_output[1822] = '{32'h305e1fe2};
/*############ DEBUG ############
test_input[14576:14583] = '{88.8490701898, 45.6913091827, 49.9831246172, -35.9057057521, 37.0471178711, -58.57587743, -97.2068253629, 67.9127156161};
test_label[1822] = '{88.8490701898};
test_output[1822] = '{8.08084377517e-10};
############ END DEBUG ############*/
test_input[14584:14591] = '{32'h429f136e, 32'h422107ce, 32'h4298e730, 32'hc287d299, 32'hc2ad95be, 32'hc28f2c0c, 32'h41f2c054, 32'hc2396297};
test_label[1823] = '{32'hc2ad95be};
test_output[1823] = '{32'h43266004};
/*############ DEBUG ############
test_input[14584:14591] = '{79.5379458708, 40.257621794, 76.4515407874, -67.9113202486, -86.7924622414, -71.5860252773, 30.3439110457, -46.3462796004};
test_label[1823] = '{-86.7924622414};
test_output[1823] = '{166.375061947};
############ END DEBUG ############*/
test_input[14592:14599] = '{32'hc2c57062, 32'hc2c1cd03, 32'hc271837b, 32'hc192bfb8, 32'hc257d2ba, 32'hc20338f7, 32'hc280ffd2, 32'hc29ff457};
test_label[1824] = '{32'hc2c57062};
test_output[1824] = '{32'h42a0c074};
/*############ DEBUG ############
test_input[14592:14599] = '{-98.7194972489, -96.9004113524, -60.378398978, -18.3436133451, -53.9557857904, -32.8056281068, -64.4996501614, -79.9772265524};
test_label[1824] = '{-98.7194972489};
test_output[1824] = '{80.3758844276};
############ END DEBUG ############*/
test_input[14600:14607] = '{32'h41963c7d, 32'hc2baea95, 32'h42107790, 32'hc224a9d8, 32'hc2946188, 32'hc160d43e, 32'hc2823475, 32'h4192ee47};
test_label[1825] = '{32'h42107790};
test_output[1825] = '{32'h3352ddf8};
/*############ DEBUG ############
test_input[14600:14607] = '{18.7795347188, -93.4581678654, 36.1167600248, -41.1658620449, -74.1904936315, -14.0518168129, -65.1024546582, 18.3663463298};
test_label[1825] = '{36.1167600248};
test_output[1825] = '{4.90963143313e-08};
############ END DEBUG ############*/
test_input[14608:14615] = '{32'hc29cbdc1, 32'hc2102c41, 32'h42000cca, 32'hc0876c50, 32'hc2107214, 32'h416dcc74, 32'hc1cb0b1a, 32'hc12ad4bf};
test_label[1826] = '{32'h416dcc74};
test_output[1826] = '{32'h4189335b};
/*############ DEBUG ############
test_input[14608:14615] = '{-78.3706162323, -36.0432175125, 32.0124909205, -4.2319719416, -36.1114048341, 14.8624148951, -25.3804214226, -10.6769400549};
test_label[1826] = '{14.8624148951};
test_output[1826] = '{17.1500760611};
############ END DEBUG ############*/
test_input[14616:14623] = '{32'hc297112b, 32'hc1d81159, 32'hc19f8fc5, 32'h427cb540, 32'h42b78e6d, 32'h42bdb227, 32'hc2870e21, 32'hc298bfad};
test_label[1827] = '{32'hc19f8fc5};
test_output[1827] = '{32'h42e5ad55};
/*############ DEBUG ############
test_input[14616:14623] = '{-75.533531485, -27.0084698556, -19.945200801, 63.1770001181, 91.7781717226, 94.8479507798, -67.5275961377, -76.3743663342};
test_label[1827] = '{-19.945200801};
test_output[1827] = '{114.838537302};
############ END DEBUG ############*/
test_input[14624:14631] = '{32'h421e3cf1, 32'hc187e510, 32'hc27eebe2, 32'hc26c89ad, 32'hc25af3ec, 32'hc29559d9, 32'h4207a09e, 32'h42b34324};
test_label[1828] = '{32'h42b34324};
test_output[1828] = '{32'h80000000};
/*############ DEBUG ############
test_input[14624:14631] = '{39.5595124134, -16.9868464526, -63.7303555681, -59.1344487457, -54.7382053973, -74.6754839624, 33.9068543619, 89.631136058};
test_label[1828] = '{89.631136058};
test_output[1828] = '{-0.0};
############ END DEBUG ############*/
test_input[14632:14639] = '{32'h4283ae13, 32'h421667a9, 32'hc21e59c9, 32'h41dc1925, 32'hc2c4d404, 32'h428fcdf2, 32'h3ec2b6d9, 32'hc2689f4c};
test_label[1829] = '{32'hc2c4d404};
test_output[1829] = '{32'h432a5194};
/*############ DEBUG ############
test_input[14632:14639] = '{65.8399924477, 37.601232392, -39.5876800324, 27.5122770121, -98.4140934918, 71.9022385093, 0.380301257924, -58.1555622125};
test_label[1829] = '{-98.4140934918};
test_output[1829] = '{170.318658456};
############ END DEBUG ############*/
test_input[14640:14647] = '{32'h425f988c, 32'hc108e859, 32'hc1babb44, 32'h42736a81, 32'h420670db, 32'hc2623613, 32'h4238749d, 32'h429b65ab};
test_label[1830] = '{32'h429b65ab};
test_output[1830] = '{32'h33512ce1};
/*############ DEBUG ############
test_input[14640:14647] = '{55.898969696, -8.55672593828, -23.3414387496, 60.8540086636, 33.6102087938, -56.5528080427, 46.1138810658, 77.6985692067};
test_label[1830] = '{77.6985692067};
test_output[1830] = '{4.87024212828e-08};
############ END DEBUG ############*/
test_input[14648:14655] = '{32'h42c43c58, 32'h41131f73, 32'hc291748a, 32'h42781942, 32'hc282db7c, 32'hc22d7832, 32'h4286c911, 32'hc2a3c98a};
test_label[1831] = '{32'h4286c911};
test_output[1831] = '{32'h41f5cd1f};
/*############ DEBUG ############
test_input[14648:14655] = '{98.1178625059, 9.19517831138, -72.7276170229, 62.0246676033, -65.4286795863, -43.3673774516, 67.3927058857, -81.8936284242};
test_label[1831] = '{67.3927058857};
test_output[1831] = '{30.7251566202};
############ END DEBUG ############*/
test_input[14656:14663] = '{32'hc2ba26f9, 32'hc2906471, 32'h42731541, 32'h42c5629c, 32'h410a8ecc, 32'h3ffffbfc, 32'h427f4361, 32'hc1b41df6};
test_label[1832] = '{32'h427f4361};
test_output[1832] = '{32'h420b81d8};
/*############ DEBUG ############
test_input[14656:14663] = '{-93.0761191754, -72.1961737096, 60.7707562566, 98.6925987565, 8.65986206695, 1.99987746681, 63.8157989575, -22.5146285624};
test_label[1832] = '{63.8157989575};
test_output[1832] = '{34.876799799};
############ END DEBUG ############*/
test_input[14664:14671] = '{32'h428cfbe3, 32'hc2a6841c, 32'h4255797d, 32'h40bc8418, 32'hc279419a, 32'h423a05cd, 32'h424ecbc5, 32'h41cdc3b7};
test_label[1833] = '{32'hc279419a};
test_output[1833] = '{32'h4304ce58};
/*############ DEBUG ############
test_input[14664:14671] = '{70.4919675909, -83.2580258654, 53.368641766, 5.89112463665, -62.3140648911, 46.5056659158, 51.698992448, 25.7205635913};
test_label[1833] = '{-62.3140648911};
test_output[1833] = '{132.806032525};
############ END DEBUG ############*/
test_input[14672:14679] = '{32'hc2257fab, 32'hc1acb10a, 32'h41e6d69f, 32'hc0119147, 32'hc25fd2ae, 32'hc192be1c, 32'hc2034e08, 32'hc26d4ef1};
test_label[1834] = '{32'hc192be1c};
test_output[1834] = '{32'h423cca5d};
/*############ DEBUG ############
test_input[14672:14679] = '{-41.3746738695, -21.5864454156, 28.8547955726, -2.2744919763, -55.955741163, -18.3428265632, -32.8262017398, -59.3270911948};
test_label[1834] = '{-18.3428265632};
test_output[1834] = '{47.1976221358};
############ END DEBUG ############*/
test_input[14680:14687] = '{32'hc2228361, 32'h420ec565, 32'h41b7cf79, 32'hc2b844f6, 32'h428d41a8, 32'h428a218d, 32'hc2865edb, 32'hc2946ee4};
test_label[1835] = '{32'hc2b844f6};
test_output[1835] = '{32'h4322f404};
/*############ DEBUG ############
test_input[14680:14687] = '{-40.6283000252, 35.6927683153, 22.976305103, -92.1346911549, 70.6282382998, 69.0655270431, -67.1852655166, -74.2165854097};
test_label[1835] = '{-92.1346911549};
test_output[1835] = '{162.95319199};
############ END DEBUG ############*/
test_input[14688:14695] = '{32'hc1a44fbb, 32'hc1e609b9, 32'hc2c030a3, 32'h42927aa4, 32'hc03221f6, 32'h42a3f030, 32'h42873ef6, 32'h4182a4ce};
test_label[1836] = '{32'hc03221f6};
test_output[1836] = '{32'h42a98155};
/*############ DEBUG ############
test_input[14688:14695] = '{-20.5389300869, -28.7547480425, -96.0949937467, 73.2395329384, -2.7833227277, 81.9691185851, 67.6229670318, 16.3304707224};
test_label[1836] = '{-2.7833227277};
test_output[1836] = '{84.7526036173};
############ END DEBUG ############*/
test_input[14696:14703] = '{32'h4208b682, 32'hc2766991, 32'hc1b73591, 32'hc2c12bc6, 32'hc13d9413, 32'hc121a044, 32'h42ab9fea, 32'hc20b165f};
test_label[1837] = '{32'hc20b165f};
test_output[1837] = '{32'h42f12b1a};
/*############ DEBUG ############
test_input[14696:14703] = '{34.1782295808, -61.6030918712, -22.901154572, -96.5854963709, -11.8486510997, -10.1016278108, 85.8123316812, -34.7718474382};
test_label[1837] = '{-34.7718474382};
test_output[1837] = '{120.584179119};
############ END DEBUG ############*/
test_input[14704:14711] = '{32'hc2b6c0d7, 32'hc29c5f91, 32'hc2c13d35, 32'h42967f4b, 32'h42b524a0, 32'h41b56718, 32'hc0c1c9a4, 32'hc1ce2243};
test_label[1838] = '{32'hc0c1c9a4};
test_output[1838] = '{32'h42c1413a};
/*############ DEBUG ############
test_input[14704:14711] = '{-91.3766415652, -78.1866554361, -96.6195449278, 75.2486195036, 90.5715320536, 22.6753383972, -6.05586453452, -25.7667291563};
test_label[1838] = '{-6.05586453452};
test_output[1838] = '{96.6273968096};
############ END DEBUG ############*/
test_input[14712:14719] = '{32'h429113da, 32'h423101fe, 32'hc139e4c2, 32'h42685c7d, 32'hc2bc4cbb, 32'h42b73c14, 32'h42bc5f58, 32'h4210790a};
test_label[1839] = '{32'h423101fe};
test_output[1839] = '{32'h4248084a};
/*############ DEBUG ############
test_input[14712:14719] = '{72.5387724514, 44.2519470441, -11.6183486883, 58.0903211636, -94.1498618392, 91.6173377819, 94.1862153107, 36.1182035338};
test_label[1839] = '{44.2519470441};
test_output[1839] = '{50.0080961666};
############ END DEBUG ############*/
test_input[14720:14727] = '{32'h42a94b20, 32'hc1387d7f, 32'h428212c5, 32'hc22e5872, 32'h429efc3a, 32'h4299a70e, 32'hc25150a5, 32'h42a3dbff};
test_label[1840] = '{32'h429efc3a};
test_output[1840] = '{32'h40a729d7};
/*############ DEBUG ############
test_input[14720:14727] = '{84.6467276557, -11.5306384655, 65.0366613468, -43.586371802, 79.4926265263, 76.8262772472, -52.3287528611, 81.9296821209};
test_label[1840] = '{79.4926265263};
test_output[1840] = '{5.22385737091};
############ END DEBUG ############*/
test_input[14728:14735] = '{32'hc2c6d741, 32'hc269bf29, 32'hc265c1a7, 32'h42929f43, 32'hc190b6d3, 32'h42b54fa1, 32'h424a7729, 32'hc281b720};
test_label[1841] = '{32'hc281b720};
test_output[1841] = '{32'h431b8360};
/*############ DEBUG ############
test_input[14728:14735] = '{-99.4204141088, -58.43668069, -57.4391125322, 73.3110597023, -18.0892700681, 90.6555262149, 50.6163690625, -64.8576638219};
test_label[1841] = '{-64.8576638219};
test_output[1841] = '{155.513190066};
############ END DEBUG ############*/
test_input[14736:14743] = '{32'hc29ced63, 32'h42b440cd, 32'h414818a3, 32'hc22de113, 32'hc16a9877, 32'hc2b58fc0, 32'h42c40a2b, 32'hc17c26ef};
test_label[1842] = '{32'h42b440cd};
test_output[1842] = '{32'h40fc98f0};
/*############ DEBUG ############
test_input[14736:14743] = '{-78.4636493053, 90.1265613327, 12.506014766, -43.469799311, -14.6622225876, -90.7807594852, 98.0198575058, -15.7595048292};
test_label[1842] = '{90.1265613327};
test_output[1842] = '{7.89366934081};
############ END DEBUG ############*/
test_input[14744:14751] = '{32'hc1faa507, 32'hc2b439cf, 32'h42b28275, 32'hc2ae3795, 32'hc189d8c6, 32'hc10ee336, 32'hc15bb5ba, 32'h42670ce9};
test_label[1843] = '{32'hc189d8c6};
test_output[1843] = '{32'h42d4f8a7};
/*############ DEBUG ############
test_input[14744:14751] = '{-31.3305797496, -90.1129049131, 89.2548020156, -87.1085577076, -17.2308468114, -8.93047122794, -13.731866954, 57.7626070269};
test_label[1843] = '{-17.2308468114};
test_output[1843] = '{106.485648827};
############ END DEBUG ############*/
test_input[14752:14759] = '{32'hbf060222, 32'h4281f559, 32'hc2b1e422, 32'h42ba504f, 32'h41fd68aa, 32'h42380672, 32'h40d60f89, 32'hc27d3548};
test_label[1844] = '{32'h40d60f89};
test_output[1844] = '{32'h42acef57};
/*############ DEBUG ############
test_input[14752:14759] = '{-0.523470044554, 64.9791950325, -88.9455751008, 93.1568534272, 31.6761062698, 46.0062933019, 6.689396271, -63.3020312587};
test_label[1844] = '{6.689396271};
test_output[1844] = '{86.4674571562};
############ END DEBUG ############*/
test_input[14760:14767] = '{32'hc2ada07e, 32'hc2aa3434, 32'hc2bb4c52, 32'hc283fdad, 32'hc2b23621, 32'h3f5144a1, 32'hc1182d1b, 32'h408d360d};
test_label[1845] = '{32'h408d360d};
test_output[1845] = '{32'h3cddd867};
/*############ DEBUG ############
test_input[14760:14767] = '{-86.8134620071, -85.1019560763, -93.6490659463, -65.9954621621, -89.1057168261, 0.817453435783, -9.51101178198, 4.41284816929};
test_label[1845] = '{4.41284816929};
test_output[1845] = '{0.0270807275311};
############ END DEBUG ############*/
test_input[14768:14775] = '{32'h42ab95a6, 32'hc27a1212, 32'hc255ca25, 32'h41b430e2, 32'h42b8ff43, 32'hc134e6f9, 32'hc274790c, 32'hc08208d3};
test_label[1846] = '{32'h42b8ff43};
test_output[1846] = '{32'h3aa03b10};
/*############ DEBUG ############
test_input[14768:14775] = '{85.7922821048, -62.5176468621, -53.4474076321, 22.5238692978, 92.4985581714, -11.3063895267, -61.1182100725, -4.0635772707};
test_label[1846] = '{92.4985581714};
test_output[1846] = '{0.00122246329635};
############ END DEBUG ############*/
test_input[14776:14783] = '{32'h42a030a8, 32'hc1906618, 32'h4129f8d4, 32'h42a6bc64, 32'h42350e4d, 32'hc20876b0, 32'hc1fe3461, 32'hc1a8b7f6};
test_label[1847] = '{32'hc1fe3461};
test_output[1847] = '{32'h42e65c87};
/*############ DEBUG ############
test_input[14776:14783] = '{80.095027994, -18.0498504037, 10.6232486571, 83.3679494866, 45.2639641195, -34.1159068552, -31.7755749315, -21.0898251949};
test_label[1847] = '{-31.7755749315};
test_output[1847] = '{115.180719575};
############ END DEBUG ############*/
test_input[14784:14791] = '{32'h418bffd5, 32'hc09c3277, 32'hc29fff64, 32'h4119d80f, 32'hc2b972ef, 32'h4297b55c, 32'hc137b6c6, 32'hbe275467};
test_label[1848] = '{32'h4297b55c};
test_output[1848] = '{32'h80000000};
/*############ DEBUG ############
test_input[14784:14791] = '{17.4999182236, -4.88116044201, -79.9988083399, 9.61524834175, -92.7244814452, 75.8542210014, -11.482122758, -0.163407905797};
test_label[1848] = '{75.8542210014};
test_output[1848] = '{-0.0};
############ END DEBUG ############*/
test_input[14792:14799] = '{32'h429b5d2c, 32'hc25f4b20, 32'h42872abe, 32'h42bc3315, 32'h42425e9b, 32'h422f539d, 32'h420298fa, 32'hc182f46e};
test_label[1849] = '{32'hc182f46e};
test_output[1849] = '{32'h42dcf031};
/*############ DEBUG ############
test_input[14792:14799] = '{77.6819784248, -55.8233650723, 67.5834829876, 94.0997718979, 48.5923871103, 43.831652217, 32.6493928592, -16.3693500972};
test_label[1849] = '{-16.3693500972};
test_output[1849] = '{110.469122069};
############ END DEBUG ############*/
test_input[14800:14807] = '{32'hc12887a4, 32'hc20f228e, 32'h421ecdde, 32'h4295d2d5, 32'h427357fb, 32'h42884172, 32'h422e5e15, 32'hc22024f2};
test_label[1850] = '{32'h42884172};
test_output[1850] = '{32'h40d91f77};
/*############ DEBUG ############
test_input[14800:14807] = '{-10.5331155683, -35.7837432409, 39.7010438473, 74.9117822962, 60.8359181521, 68.1278234969, 43.5918773339, -40.0360777177};
test_label[1850] = '{68.1278234969};
test_output[1850] = '{6.78509071469};
############ END DEBUG ############*/
test_input[14808:14815] = '{32'h42861ba0, 32'hc2018346, 32'hc1b1f109, 32'hc2be04a4, 32'h41bea5bb, 32'hc2320481, 32'h40848604, 32'h40930bd3};
test_label[1851] = '{32'h41bea5bb};
test_output[1851] = '{32'h422ce462};
/*############ DEBUG ############
test_input[14808:14815] = '{67.0539516163, -32.3781983324, -22.2426933653, -95.0090624323, 23.8309222847, -44.504398256, 4.14135952737, 4.59519323446};
test_label[1851] = '{23.8309222847};
test_output[1851] = '{43.2230293317};
############ END DEBUG ############*/
test_input[14816:14823] = '{32'h41e734b9, 32'h41f6d6c7, 32'h42b55324, 32'h42afb6fb, 32'hc20fbf7c, 32'hc2827fc0, 32'h42a8e27a, 32'hc29dbf9d};
test_label[1852] = '{32'h42a8e27a};
test_output[1852] = '{32'h40c8fb36};
/*############ DEBUG ############
test_input[14816:14823] = '{28.9007426396, 30.8548725187, 90.6623824909, 87.8573812065, -35.9369957225, -65.2495117334, 84.4423379952, -78.8742471851};
test_label[1852] = '{84.4423379952};
test_output[1852] = '{6.28066521176};
############ END DEBUG ############*/
test_input[14824:14831] = '{32'h4251ec16, 32'hc2379561, 32'h42c428b4, 32'h429a63b9, 32'h428dcf2f, 32'h422b0bb8, 32'hc2c2610a, 32'h42708711};
test_label[1853] = '{32'h422b0bb8};
test_output[1853] = '{32'h425d45b0};
/*############ DEBUG ############
test_input[14824:14831] = '{52.4805544625, -45.8958791121, 98.0795012989, 77.1947685591, 70.904656101, 42.7614452331, -97.1895313973, 60.1319000546};
test_label[1853] = '{42.7614452331};
test_output[1853] = '{55.3180560667};
############ END DEBUG ############*/
test_input[14832:14839] = '{32'hc1662473, 32'hc03f434c, 32'h427df696, 32'h418c855d, 32'hc0e6a464, 32'h42388808, 32'hc284659b, 32'hc206e2ba};
test_label[1854] = '{32'h427df696};
test_output[1854] = '{32'h32f89c85};
/*############ DEBUG ############
test_input[14832:14839] = '{-14.3838984692, -2.98848249337, 63.4908078681, 17.5651188198, -7.20756734385, 46.132841999, -66.1984506989, -33.7214117842};
test_label[1854] = '{63.4908078681};
test_output[1854] = '{2.89421772961e-08};
############ END DEBUG ############*/
test_input[14840:14847] = '{32'hc2b2ad2e, 32'hc12ae676, 32'hc253efda, 32'hc2b60e31, 32'h42197bdc, 32'hbf74e85f, 32'h42269dd8, 32'h423a18dc};
test_label[1855] = '{32'hc12ae676};
test_output[1855] = '{32'h4264da98};
/*############ DEBUG ############
test_input[14840:14847] = '{-89.3382427963, -10.6812651434, -52.9842300248, -91.0277159709, 38.3709558091, -0.956670676828, 41.654144855, 46.5242775833};
test_label[1855] = '{-10.6812651434};
test_output[1855] = '{57.2134713367};
############ END DEBUG ############*/
test_input[14848:14855] = '{32'h41dca574, 32'hc1ec25dd, 32'hc2c1df3f, 32'h413eda1e, 32'hc2bb997e, 32'hc2bc9a46, 32'hc19b73a6, 32'h429b7f65};
test_label[1856] = '{32'h413eda1e};
test_output[1856] = '{32'h4283a421};
/*############ DEBUG ############
test_input[14848:14855] = '{27.5807867582, -29.5184883305, -96.9360284978, 11.9282511581, -93.7997920974, -94.3013160087, -19.4314693901, 77.7488158316};
test_label[1856] = '{11.9282511581};
test_output[1856] = '{65.8205646735};
############ END DEBUG ############*/
test_input[14856:14863] = '{32'h3f8fe319, 32'hc197dfff, 32'h42c06ca3, 32'h42c098dc, 32'h41d8a76d, 32'h42859ee9, 32'hc2546cee, 32'h418f7553};
test_label[1857] = '{32'h42859ee9};
test_output[1857] = '{32'h41f11cd3};
/*############ DEBUG ############
test_input[14856:14863] = '{1.12411791292, -18.984373505, 96.2121842031, 96.2985520879, 27.0817517133, 66.8103727959, -53.1063749968, 17.9322881214};
test_label[1857] = '{66.8103727959};
test_output[1857] = '{30.1390746669};
############ END DEBUG ############*/
test_input[14864:14871] = '{32'h419890c0, 32'hc2622880, 32'hc0fdae12, 32'h428c8576, 32'hc29e09e1, 32'h421e5a95, 32'hc2aa317e, 32'hc24b6414};
test_label[1858] = '{32'h428c8576};
test_output[1858] = '{32'h29570000};
/*############ DEBUG ############
test_input[14864:14871] = '{19.0706796267, -56.5395505822, -7.92749870438, 70.2606677911, -79.0192968507, 39.5884607826, -85.0966625797, -50.8477337992};
test_label[1858] = '{70.2606677911};
test_output[1858] = '{4.77395900589e-14};
############ END DEBUG ############*/
test_input[14872:14879] = '{32'hc26cae26, 32'h42830f65, 32'h40e6c9a6, 32'h414d2ee5, 32'hc22946e4, 32'h3f0d8632, 32'h421cf624, 32'hc29c9041};
test_label[1859] = '{32'h42830f65};
test_output[1859] = '{32'h2c868d00};
/*############ DEBUG ############
test_input[14872:14879] = '{-59.1700687352, 65.5300661103, 7.21211538127, 12.8239492138, -42.3192288514, 0.552828923256, 39.2403700901, -78.2817487435};
test_label[1859] = '{65.5300661103};
test_output[1859] = '{3.82416320833e-12};
############ END DEBUG ############*/
test_input[14880:14887] = '{32'h42a448ac, 32'hc29d49a2, 32'h424136a5, 32'hc186dbb0, 32'hc2b048ff, 32'h429418e9, 32'hc1e7ec0c, 32'hc147d086};
test_label[1860] = '{32'h42a448ac};
test_output[1860] = '{32'h39a03092};
/*############ DEBUG ############
test_input[14880:14887] = '{82.1419383618, -78.6438170844, 48.3033630827, -16.8572686746, -88.1425675672, 74.0486535769, -28.9902576719, -12.488408726};
test_label[1860] = '{82.1419383618};
test_output[1860] = '{0.000305537646568};
############ END DEBUG ############*/
test_input[14888:14895] = '{32'h410dcd87, 32'h42437c1f, 32'h41eca51c, 32'hc11d0908, 32'h3f69d7a6, 32'hc292183c, 32'hc2ab211e, 32'h41aaacec};
test_label[1861] = '{32'hc292183c};
test_output[1861] = '{32'h42f3d64b};
/*############ DEBUG ############
test_input[14888:14895] = '{8.86267772791, 48.8712127512, 29.5806189682, -9.81470492711, 0.913446774755, -73.0473313575, -85.5646839678, 21.3344347777};
test_label[1861] = '{-73.0473313575};
test_output[1861] = '{121.918544113};
############ END DEBUG ############*/
test_input[14896:14903] = '{32'h41c7d1b8, 32'hc1bbf6f5, 32'hc2b0025c, 32'hc2815be5, 32'hc2296a21, 32'h423968e0, 32'h42a5eb47, 32'h426c4f47};
test_label[1862] = '{32'hc2296a21};
test_output[1862] = '{32'h42faa058};
/*############ DEBUG ############
test_input[14896:14903] = '{24.9774022859, -23.4955840062, -88.0046103024, -64.6794851963, -42.3536403214, 46.352415515, 82.9595292706, 59.0774177439};
test_label[1862] = '{-42.3536403214};
test_output[1862] = '{125.313169592};
############ END DEBUG ############*/
test_input[14904:14911] = '{32'h42a6c12d, 32'h421231b2, 32'h422d0b96, 32'h41205b66, 32'hc1ab153e, 32'h4208e461, 32'hc219db68, 32'hc2669983};
test_label[1863] = '{32'h421231b2};
test_output[1863] = '{32'h423b50a8};
/*############ DEBUG ############
test_input[14904:14911] = '{83.3772945423, 36.5485304716, 43.2613130992, 10.0223139003, -21.385371257, 34.2230276315, -38.4642620372, -57.6499145639};
test_label[1863] = '{36.5485304716};
test_output[1863] = '{46.8287640707};
############ END DEBUG ############*/
test_input[14912:14919] = '{32'hc2a469e3, 32'h4148b5c3, 32'h42a6f6fc, 32'h429d3955, 32'hc297a67a, 32'h42514248, 32'hc1c5276d, 32'hc0f29b42};
test_label[1864] = '{32'hc2a469e3};
test_output[1864] = '{32'h4325b264};
/*############ DEBUG ############
test_input[14912:14919] = '{-82.2068095387, 12.5443751165, 83.4823888378, 78.6119740487, -75.8251499997, 52.3147267106, -24.6442517027, -7.58145238233};
test_label[1864] = '{-82.2068095387};
test_output[1864] = '{165.696839293};
############ END DEBUG ############*/
test_input[14920:14927] = '{32'h406ec549, 32'h41d8fb75, 32'hc289d066, 32'hc175f437, 32'h40bff474, 32'h428e7fae, 32'h422ba504, 32'hc172af2e};
test_label[1865] = '{32'h428e7fae};
test_output[1865] = '{32'h2b0ac800};
/*############ DEBUG ############
test_input[14920:14927] = '{3.73079142159, 27.1227816718, -68.907024568, -15.3721230538, 5.99859043494, 71.2493730871, 42.9111471996, -15.1677683211};
test_label[1865] = '{71.2493730871};
test_output[1865] = '{4.93050045236e-13};
############ END DEBUG ############*/
test_input[14928:14935] = '{32'h42584756, 32'h42bb5425, 32'hc2c7456b, 32'h428f28ac, 32'h413fd8bc, 32'h42912ee4, 32'h429ce281, 32'hc26380d9};
test_label[1866] = '{32'hc26380d9};
test_output[1866] = '{32'h43168a49};
/*############ DEBUG ############
test_input[14928:14935] = '{54.0696637739, 93.6643464027, -99.6355845243, 71.5794374234, 11.9904133373, 72.5915856557, 78.4423907907, -56.8758290072};
test_label[1866] = '{-56.8758290072};
test_output[1866] = '{150.540175656};
############ END DEBUG ############*/
test_input[14936:14943] = '{32'hc24bf23e, 32'h42424a84, 32'hc1b655ef, 32'h42bb7652, 32'hc2a3151a, 32'hc28ed930, 32'h418a1775, 32'hc1fe7488};
test_label[1867] = '{32'hc2a3151a};
test_output[1867] = '{32'h432f45b6};
/*############ DEBUG ############
test_input[14936:14943] = '{-50.9865638293, 48.5727692903, -22.7919595138, 93.7310934164, -81.5412150498, -71.4241963713, 17.2614534943, -31.806899729};
test_label[1867] = '{-81.5412150498};
test_output[1867] = '{175.272308466};
############ END DEBUG ############*/
test_input[14944:14951] = '{32'h42be689d, 32'hc1b51860, 32'h428e7626, 32'h4030f0d3, 32'hc195448a, 32'hc2723b8a, 32'h421f3352, 32'hc1d7c692};
test_label[1868] = '{32'h42be689d};
test_output[1868] = '{32'h2e2a7b20};
/*############ DEBUG ############
test_input[14944:14951] = '{95.2043214519, -22.636900905, 71.2307620186, 2.76469864698, -18.6584665503, -60.5581447535, 39.8001156334, -26.9719580349};
test_label[1868] = '{95.2043214519};
test_output[1868] = '{3.8762881794e-11};
############ END DEBUG ############*/
test_input[14952:14959] = '{32'h41f481fd, 32'h42289139, 32'hc28d002a, 32'h4298072f, 32'hc2adb08d, 32'h4153b454, 32'hc250a6b8, 32'h410fb61d};
test_label[1869] = '{32'h41f481fd};
test_output[1869] = '{32'h4235cd5f};
/*############ DEBUG ############
test_input[14952:14959] = '{30.5634716678, 42.1418195026, -70.5003197269, 76.0140299256, -86.84482952, 13.231525517, -52.1628100781, 8.98196159691};
test_label[1869] = '{30.5634716678};
test_output[1869] = '{45.4505582578};
############ END DEBUG ############*/
test_input[14960:14967] = '{32'h41752b2d, 32'h426edc60, 32'h42c3f59a, 32'hc2b4b60c, 32'hc242f768, 32'hc2c21c4c, 32'hc280f91e, 32'h428f7f5a};
test_label[1870] = '{32'h428f7f5a};
test_output[1870] = '{32'h41d1d900};
/*############ DEBUG ############
test_input[14960:14967] = '{15.3230413028, 59.7152086851, 97.9796891783, -90.3555585109, -48.7416065464, -97.0552711345, -64.4865582304, 71.748732444};
test_label[1870] = '{71.748732444};
test_output[1870] = '{26.2309567343};
############ END DEBUG ############*/
test_input[14968:14975] = '{32'hc2a73f00, 32'hc2ad3e94, 32'hc2badafa, 32'h41eab9a6, 32'h428a3de3, 32'hc1cadef6, 32'hc24d7e09, 32'hc20cd81f};
test_label[1871] = '{32'hc2badafa};
test_output[1871] = '{32'h43228c6f};
/*############ DEBUG ############
test_input[14968:14975] = '{-83.6230437398, -86.6222192422, -93.4276923178, 29.3406491417, 69.1208743712, -25.3588669284, -51.3730821625, -35.2110569822};
test_label[1871] = '{-93.4276923178};
test_output[1871] = '{162.548566689};
############ END DEBUG ############*/
test_input[14976:14983] = '{32'h4220bbe1, 32'h42bab965, 32'hc29e4014, 32'h4183851b, 32'h4272e2de, 32'hc273c49c, 32'hc21680ff, 32'h41a48c31};
test_label[1872] = '{32'h41a48c31};
test_output[1872] = '{32'h42919659};
/*############ DEBUG ############
test_input[14976:14983] = '{40.1834765331, 93.3621005247, -79.1251508751, 16.4399936409, 60.7215492928, -60.9420015512, -37.625972916, 20.5684524381};
test_label[1872] = '{20.5684524381};
test_output[1872] = '{72.7936480866};
############ END DEBUG ############*/
test_input[14984:14991] = '{32'hc1e8ce76, 32'hc2af8e8f, 32'hc27d2b46, 32'h406eaf62, 32'hc25fa6ac, 32'h4218533e, 32'h427b43b0, 32'h42674246};
test_label[1873] = '{32'h42674246};
test_output[1873] = '{32'h40a0423c};
/*############ DEBUG ############
test_input[14984:14991] = '{-29.1008106489, -87.7784326973, -63.2922576962, 3.72945449554, -55.9127662091, 38.0812895338, 62.8161008778, 57.8147219376};
test_label[1873] = '{57.8147219376};
test_output[1873] = '{5.00808506605};
############ END DEBUG ############*/
test_input[14992:14999] = '{32'hc2b843e2, 32'hc277ae62, 32'h4259e3e4, 32'h42887e4e, 32'hc23d32b4, 32'hc2a7fce1, 32'hc12e5040, 32'hc190ebeb};
test_label[1874] = '{32'hc2b843e2};
test_output[1874] = '{32'h43206118};
/*############ DEBUG ############
test_input[14992:14999] = '{-92.1325810433, -61.9202955596, 54.4725478041, 68.2466885354, -47.2995166372, -83.993902445, -10.8945922187, -18.1151939328};
test_label[1874] = '{-92.1325810433};
test_output[1874] = '{160.379270621};
############ END DEBUG ############*/
test_input[15000:15007] = '{32'h4260f9b5, 32'hc1d88f1b, 32'hc2bd2ab3, 32'h42bb1d69, 32'hc1c0697b, 32'h4299e32e, 32'hc2946533, 32'h42b4fddc};
test_label[1875] = '{32'h42b4fddc};
test_output[1875] = '{32'h4046df1e};
/*############ DEBUG ############
test_input[15000:15007] = '{56.2438527241, -27.069875714, -94.5833944927, 93.5574401447, -24.0515042096, 76.9437070613, -74.1976566283, 90.4958214199};
test_label[1875] = '{90.4958214199};
test_output[1875] = '{3.10736800278};
############ END DEBUG ############*/
test_input[15008:15015] = '{32'hc2c18e75, 32'h40892581, 32'hc2bd0557, 32'hc21f040a, 32'hc29d65c1, 32'h40750ef9, 32'hc203316d, 32'h4258bd28};
test_label[1876] = '{32'hc2c18e75};
test_output[1876] = '{32'h4316f684};
/*############ DEBUG ############
test_input[15008:15015] = '{-96.7782376083, 4.28582805796, -94.5104280007, -39.7539444078, -78.6987382293, 3.82903881421, -32.7982664003, 54.1847211432};
test_label[1876] = '{-96.7782376083};
test_output[1876] = '{150.962958751};
############ END DEBUG ############*/
test_input[15016:15023] = '{32'hc1280670, 32'h429dab83, 32'h4240e2e1, 32'hc242a1ce, 32'hc26f4d9c, 32'hc239fc4a, 32'h3faa2bd3, 32'h420700f0};
test_label[1877] = '{32'h429dab83};
test_output[1877] = '{32'h29648000};
/*############ DEBUG ############
test_input[15016:15023] = '{-10.5015712364, 78.8349845552, 48.2215611741, -48.6580126755, -59.8257898642, -46.496374588, 1.32946246414, 33.7509145982};
test_label[1877] = '{78.8349845552};
test_output[1877] = '{5.07371922254e-14};
############ END DEBUG ############*/
test_input[15024:15031] = '{32'hc24405c5, 32'h423af6c1, 32'hc28270a6, 32'h42551e2c, 32'hc07b08c3, 32'hc1064b6c, 32'h4293a850, 32'hc28478f9};
test_label[1878] = '{32'hc24405c5};
test_output[1878] = '{32'h42f5ab33};
/*############ DEBUG ############
test_input[15024:15031] = '{-49.0056349273, 46.7409698367, -65.2200196722, 53.2794648419, -3.92240967586, -8.39341311264, 73.8287369348, -66.2362714542};
test_label[1878] = '{-49.0056349273};
test_output[1878] = '{122.834371863};
############ END DEBUG ############*/
test_input[15032:15039] = '{32'hc294fcd5, 32'hc1a37ae8, 32'h4194c132, 32'h42b8f7b6, 32'h42b768c3, 32'hc26ff506, 32'hc2b36b70, 32'hc271dd76};
test_label[1879] = '{32'hc271dd76};
test_output[1879] = '{32'h431953e3};
/*############ DEBUG ############
test_input[15032:15039] = '{-74.4938156238, -20.435012312, 18.5943327289, 92.4838099235, 91.7046156648, -59.9892808358, -89.7098354447, -60.4662706647};
test_label[1879] = '{-60.4662706647};
test_output[1879] = '{153.327677985};
############ END DEBUG ############*/
test_input[15040:15047] = '{32'hc12208f9, 32'h42a0560f, 32'hc19328cc, 32'hc2b89755, 32'h418fd6be, 32'hc23e0de6, 32'hc17f1eaf, 32'hc2918b2b};
test_label[1880] = '{32'hc17f1eaf};
test_output[1880] = '{32'h42c039e5};
/*############ DEBUG ############
test_input[15040:15047] = '{-10.1271903106, 80.1680844904, -18.3949198791, -92.2955720878, 17.979855338, -47.513572032, -15.9449911145, -72.7718134117};
test_label[1880] = '{-15.9449911145};
test_output[1880] = '{96.1130756049};
############ END DEBUG ############*/
test_input[15048:15055] = '{32'h4298a7c6, 32'h408665f5, 32'hc1c9dcbc, 32'hc2b80cd6, 32'h42182d36, 32'hc2983ccd, 32'hc2a97545, 32'hc1fb2faf};
test_label[1881] = '{32'h408665f5};
test_output[1881] = '{32'h42904167};
/*############ DEBUG ############
test_input[15048:15055] = '{76.3276844003, 4.19994601248, -25.2327809162, -92.0250715745, 38.0441532082, -76.1187548548, -84.7290408417, -31.3982828063};
test_label[1881] = '{4.19994601248};
test_output[1881] = '{72.1277383878};
############ END DEBUG ############*/
test_input[15056:15063] = '{32'hc1dec0be, 32'h405a5016, 32'h41801f2a, 32'h429d602a, 32'h4242b2de, 32'h40ae6f8d, 32'hc2c5722c, 32'hbfbd6ddb};
test_label[1882] = '{32'hc2c5722c};
test_output[1882] = '{32'h4331692b};
/*############ DEBUG ############
test_input[15056:15063] = '{-27.8441120322, 3.41113799003, 16.0152171113, 78.6878204032, 48.6746763354, 5.45111714879, -98.7229949838, -1.47991502966};
test_label[1882] = '{-98.7229949838};
test_output[1882] = '{177.410815387};
############ END DEBUG ############*/
test_input[15064:15071] = '{32'h41bd8327, 32'hc28f2e56, 32'hc2c340d1, 32'hc1ea632d, 32'h41e8cb61, 32'hc2411225, 32'h421e5078, 32'h41b6dc8c};
test_label[1883] = '{32'h41bd8327};
test_output[1883] = '{32'h417e3baf};
/*############ DEBUG ############
test_input[15064:15071] = '{23.6890400507, -71.5904976698, -97.6265937165, -29.2984257952, 29.0993052187, -48.2677192624, 39.5785831195, 22.8576887036};
test_label[1883] = '{23.6890400507};
test_output[1883] = '{15.8895713618};
############ END DEBUG ############*/
test_input[15072:15079] = '{32'h4103844f, 32'h42bb0b68, 32'hc0ecbc5b, 32'hc2b16ef7, 32'h423d3007, 32'h428968cc, 32'h428563f8, 32'hc1df44f3};
test_label[1884] = '{32'h42bb0b68};
test_output[1884] = '{32'h2da64200};
/*############ DEBUG ############
test_input[15072:15079] = '{8.21980221683, 93.5222794614, -7.39799278135, -88.7167285753, 47.2969028941, 68.7046792463, 66.6952541549, -27.9086672175};
test_label[1884] = '{93.5222794614};
test_output[1884] = '{1.89013249498e-11};
############ END DEBUG ############*/
test_input[15080:15087] = '{32'hc29ebc88, 32'h428b0299, 32'h42829a26, 32'h42987280, 32'h42b36aa4, 32'h41f21868, 32'h41c7731f, 32'hc25d57d8};
test_label[1885] = '{32'h41c7731f};
test_output[1885] = '{32'h42818ddd};
/*############ DEBUG ############
test_input[15080:15087] = '{-79.3682272347, 69.5050718549, 65.3010692556, 76.2236305561, 89.7082854484, 30.2619161683, 24.9312112373, -55.3357850808};
test_label[1885] = '{24.9312112373};
test_output[1885] = '{64.7770756049};
############ END DEBUG ############*/
test_input[15088:15095] = '{32'hc268c214, 32'hc27cb0c7, 32'hc2a3d325, 32'h427dbea1, 32'hc218ebaf, 32'h4011b1e4, 32'h4286ec21, 32'h41f93342};
test_label[1886] = '{32'h427dbea1};
test_output[1886] = '{32'h40815e16};
/*############ DEBUG ############
test_input[15088:15095] = '{-58.1895311077, -63.1726327772, -81.9123902679, 63.4361627284, -38.2301604363, 2.27648248346, 67.4611927301, 31.1500288609};
test_label[1886] = '{63.4361627284};
test_output[1886] = '{4.04273522332};
############ END DEBUG ############*/
test_input[15096:15103] = '{32'h42c0571d, 32'hc2bf1a08, 32'h40c87868, 32'hc2163584, 32'hc2646b96, 32'hc28c8dfb, 32'h4223f73a, 32'hc28560e7};
test_label[1887] = '{32'h42c0571d};
test_output[1887] = '{32'h80000000};
/*############ DEBUG ############
test_input[15096:15103] = '{96.1701445176, -95.5508389983, 6.2646980486, -37.5522616233, -57.1050637269, -70.277307978, 40.991431948, -66.6892638971};
test_label[1887] = '{96.1701445176};
test_output[1887] = '{-0.0};
############ END DEBUG ############*/
test_input[15104:15111] = '{32'hc034ccf8, 32'hc2a44a8a, 32'h41e20cb2, 32'h42c3775b, 32'hc1624ed8, 32'hc2b7caff, 32'hc257ff6b, 32'hba56ca2e};
test_label[1888] = '{32'hc2a44a8a};
test_output[1888] = '{32'h4333e0f3};
/*############ DEBUG ############
test_input[15104:15111] = '{-2.82501040196, -82.1455875031, 28.2561981386, 97.7331149465, -14.1442492044, -91.8964769175, -53.9994333246, -0.000819357909521};
test_label[1888] = '{-82.1455875031};
test_output[1888] = '{179.87870245};
############ END DEBUG ############*/
test_input[15112:15119] = '{32'hc27387c6, 32'h40b7bb2a, 32'h419df741, 32'hc2b29d52, 32'h428d5ab8, 32'h422755b2, 32'hc26de0dc, 32'hc19e4974};
test_label[1889] = '{32'hc2b29d52};
test_output[1889] = '{32'h431ffc05};
/*############ DEBUG ############
test_input[15112:15119] = '{-60.8825910819, 5.74159713501, 19.7457290522, -89.3072643441, 70.6771835985, 41.833685758, -59.4695901619, -19.7858654187};
test_label[1889] = '{-89.3072643441};
test_output[1889] = '{159.984447943};
############ END DEBUG ############*/
test_input[15120:15127] = '{32'h41833724, 32'hc2a88b9b, 32'hc2b5479d, 32'h416e2d8d, 32'h420cc3ab, 32'h42154136, 32'h424aeeff, 32'h41a98e86};
test_label[1890] = '{32'h416e2d8d};
test_output[1890] = '{32'h420f639c};
/*############ DEBUG ############
test_input[15120:15127] = '{16.4019246159, -84.2726657385, -90.6398697483, 14.8861211898, 35.1910802048, 37.3136831553, 50.7333928705, 21.1945912081};
test_label[1890] = '{14.8861211898};
test_output[1890] = '{35.8472733441};
############ END DEBUG ############*/
test_input[15128:15135] = '{32'h40a6ea9e, 32'h42819016, 32'hc20fe92e, 32'h426e5b8d, 32'hc26c6b78, 32'hc1a7de25, 32'hc2b7a00c, 32'h42a34dfe};
test_label[1891] = '{32'h42819016};
test_output[1891] = '{32'h4186f7a2};
/*############ DEBUG ############
test_input[15128:15135] = '{5.21613963011, 64.7814155281, -35.9777147013, 59.5894060898, -59.1049503173, -20.9834682758, -91.8125906417, 81.652329923};
test_label[1891] = '{64.7814155281};
test_output[1891] = '{16.8709144423};
############ END DEBUG ############*/
test_input[15136:15143] = '{32'h42b37239, 32'h4225337b, 32'h41e1875e, 32'h4198c2c1, 32'h405d7f7a, 32'h3fe3a137, 32'h4270ac32, 32'h427d0400};
test_label[1892] = '{32'h4198c2c1};
test_output[1892] = '{32'h428d4188};
/*############ DEBUG ############
test_input[15136:15143] = '{89.7230895132, 41.3002721723, 28.1910974783, 19.0950952599, 3.46090565793, 1.7783573698, 60.1681594984, 63.2539046172};
test_label[1892] = '{19.0950952599};
test_output[1892] = '{70.6279942533};
############ END DEBUG ############*/
test_input[15144:15151] = '{32'h42b2999d, 32'hc0d2db32, 32'h427d3144, 32'h4132958e, 32'h428d9490, 32'h424b989e, 32'h42ae4ce7, 32'h3fb26a54};
test_label[1893] = '{32'h42ae4ce7};
test_output[1893] = '{32'h4010a44e};
/*############ DEBUG ############
test_input[15144:15151] = '{89.3000256056, -6.58925705011, 63.298111655, 11.1615127599, 70.7901637848, 50.8990410937, 87.1501999253, 1.39386983007};
test_label[1893] = '{87.1501999253};
test_output[1893] = '{2.26002847992};
############ END DEBUG ############*/
test_input[15152:15159] = '{32'hc2a5e8c5, 32'hc298816b, 32'hc190f6ae, 32'h420fa308, 32'h422bc652, 32'h42a4892d, 32'hc10652f5, 32'h42968f11};
test_label[1894] = '{32'h422bc652};
test_output[1894] = '{32'h421d4cf9};
/*############ DEBUG ############
test_input[15152:15159] = '{-82.9546248346, -76.2527671779, -18.1204486151, 35.9092119566, 42.9436725392, 82.2679208366, -8.39525325793, 75.2794266136};
test_label[1894] = '{42.9436725392};
test_output[1894] = '{39.3251703066};
############ END DEBUG ############*/
test_input[15160:15167] = '{32'hc20f2309, 32'h423b81db, 32'hc291255e, 32'h429a3622, 32'hc14c1da0, 32'h42975f18, 32'h427b0629, 32'h4123ca24};
test_label[1895] = '{32'h4123ca24};
test_output[1895] = '{32'h42862bb6};
/*############ DEBUG ############
test_input[15160:15167] = '{-35.7842156909, 46.8768138379, -72.5729800901, 77.1057314458, -12.7572328855, 75.6857290547, 62.7560158783, 10.2368512083};
test_label[1895] = '{10.2368512083};
test_output[1895] = '{67.085372941};
############ END DEBUG ############*/
test_input[15168:15175] = '{32'hc1424076, 32'hc1efd135, 32'h424a1de8, 32'h42a7ae05, 32'h4217a411, 32'h42181cc5, 32'hc2b0c718, 32'h425279b8};
test_label[1896] = '{32'h424a1de8};
test_output[1896] = '{32'h42053e21};
/*############ DEBUG ############
test_input[15168:15175] = '{-12.1407375715, -29.9771518811, 50.5292049884, 83.8398788543, 37.9102194501, 38.0280937556, -88.3888556399, 52.6188648936};
test_label[1896] = '{50.5292049884};
test_output[1896] = '{33.3106738659};
############ END DEBUG ############*/
test_input[15176:15183] = '{32'hc281cbcf, 32'h4185281f, 32'hc2bc423c, 32'h42a1fec4, 32'h41649707, 32'hc23b116c, 32'h4279f916, 32'hc2aa2762};
test_label[1897] = '{32'h42a1fec4};
test_output[1897] = '{32'h321e02d9};
/*############ DEBUG ############
test_input[15176:15183] = '{-64.8980669189, 16.6445903241, -94.1293612349, 80.9975874626, 14.2868720276, -46.7670135367, 62.4932487735, -85.0769195484};
test_label[1897] = '{80.9975874626};
test_output[1897] = '{9.19745794869e-09};
############ END DEBUG ############*/
test_input[15184:15191] = '{32'h42bad289, 32'h42946a3f, 32'h40efe8f7, 32'hc2967903, 32'h42c35186, 32'hc29a71dd, 32'hc283d2c4, 32'h4225b1f8};
test_label[1898] = '{32'hc2967903};
test_output[1898] = '{32'h432ce8e7};
/*############ DEBUG ############
test_input[15184:15191] = '{93.4111982859, 74.2075142882, 7.49718813763, -75.2363511089, 97.6592287009, -77.2223891987, -65.9116498109, 41.4237959721};
test_label[1898] = '{-75.2363511089};
test_output[1898] = '{172.909770993};
############ END DEBUG ############*/
test_input[15192:15199] = '{32'hc22df66d, 32'h424fe7d1, 32'hc2c32440, 32'hc1dee11a, 32'hc1a483f1, 32'h42c162fc, 32'hc12e5156, 32'hc2472104};
test_label[1899] = '{32'hc2472104};
test_output[1899] = '{32'h431279bf};
/*############ DEBUG ############
test_input[15192:15199] = '{-43.4906497373, 51.9763826596, -97.5708027967, -27.8599127986, -20.5644244306, 96.6933313223, -10.8948577214, -49.7822407009};
test_label[1899] = '{-49.7822407009};
test_output[1899] = '{146.475572023};
############ END DEBUG ############*/
test_input[15200:15207] = '{32'hc28cc5b2, 32'hbe8697c4, 32'h427cf5a2, 32'hc231a90c, 32'h420e9725, 32'hc19f2d6e, 32'h424cd2f7, 32'hc2505a46};
test_label[1900] = '{32'h424cd2f7};
test_output[1900] = '{32'h41408ab0};
/*############ DEBUG ############
test_input[15200:15207] = '{-70.386121425, -0.262876631824, 63.2398743521, -44.415085982, 35.6476005783, -19.8971828111, 51.206020854, -52.0881593566};
test_label[1900] = '{51.206020854};
test_output[1900] = '{12.0338594377};
############ END DEBUG ############*/
test_input[15208:15215] = '{32'hc292fc49, 32'hc27ad849, 32'h41410cf0, 32'hc28538bb, 32'h4263b789, 32'hc2a71e1f, 32'h42a9e1fd, 32'h4225d761};
test_label[1901] = '{32'hc292fc49};
test_output[1901] = '{32'h431e6f23};
/*############ DEBUG ############
test_input[15208:15215] = '{-73.4927447954, -62.7112146748, 12.0656588457, -66.6108019421, 56.9292325369, -83.5588279818, 84.9413830402, 41.460332723};
test_label[1901] = '{-73.4927447954};
test_output[1901] = '{158.434127836};
############ END DEBUG ############*/
test_input[15216:15223] = '{32'hc24fb786, 32'hc2682781, 32'hc27b5287, 32'h42538b13, 32'h416ce0b4, 32'h427140b4, 32'h4299da6b, 32'hc1f089e9};
test_label[1902] = '{32'h4299da6b};
test_output[1902] = '{32'h3382f0e0};
/*############ DEBUG ############
test_input[15216:15223] = '{-51.9292216859, -58.0385772072, -62.8305915622, 52.8858135481, 14.8048587512, 60.3131867331, 76.9265976327, -30.0673385818};
test_label[1902] = '{76.9265976327};
test_output[1902] = '{6.09741179484e-08};
############ END DEBUG ############*/
test_input[15224:15231] = '{32'h426d6f48, 32'hc19a3040, 32'hc2afb022, 32'h421683ef, 32'h41b57d03, 32'h4183bfb8, 32'h4163fd2d, 32'h428d5599};
test_label[1903] = '{32'h4183bfb8};
test_output[1903] = '{32'h4258cb58};
/*############ DEBUG ############
test_input[15224:15231] = '{59.3586734413, -19.2735600192, -87.8440058209, 37.6288421836, 22.6860413864, 16.4686133546, 14.249310663, 70.6671805229};
test_label[1903] = '{16.4686133546};
test_output[1903] = '{54.1985794363};
############ END DEBUG ############*/
test_input[15232:15239] = '{32'h42aa8a23, 32'h4270ecdc, 32'hc1f1ff2e, 32'hc22cc6c2, 32'hc2a47f59, 32'h41089bbc, 32'h41485862, 32'hc13260a4};
test_label[1904] = '{32'h41485862};
test_output[1904] = '{32'h42917f17};
/*############ DEBUG ############
test_input[15232:15239] = '{85.2698008207, 60.2313074544, -30.249600208, -43.1941000872, -82.2487262264, 8.53802097694, 12.5215774671, -11.14859425};
test_label[1904] = '{12.5215774671};
test_output[1904] = '{72.7482233536};
############ END DEBUG ############*/
test_input[15240:15247] = '{32'hc2b12e4d, 32'h42617cbe, 32'h41834627, 32'h428ab09d, 32'h426f3f8b, 32'h4290f2f5, 32'hc25d04f6, 32'hc29778d5};
test_label[1905] = '{32'h428ab09d};
test_output[1905] = '{32'h404b0871};
/*############ DEBUG ############
test_input[15240:15247] = '{-88.5904300655, 56.3718181397, 16.4092543924, 69.3449469019, 59.8120521599, 72.4745271891, -55.2548432031, -75.7360009227};
test_label[1905] = '{69.3449469019};
test_output[1905] = '{3.17239014724};
############ END DEBUG ############*/
test_input[15248:15255] = '{32'h425eea9e, 32'h42b95342, 32'h42aa953f, 32'hc2972a5a, 32'hc21a06d7, 32'hc266470f, 32'h423f6222, 32'h4277e04b};
test_label[1906] = '{32'h4277e04b};
test_output[1906] = '{32'h41f58dbd};
/*############ DEBUG ############
test_input[15248:15255] = '{55.7291187146, 92.6626157894, 85.2914977344, -75.5827212553, -38.5066789814, -57.569391338, 47.845831447, 61.9690363485};
test_label[1906] = '{61.9690363485};
test_output[1906] = '{30.6942084073};
############ END DEBUG ############*/
test_input[15256:15263] = '{32'h4192a38a, 32'hc20ce309, 32'h429b02e2, 32'hc2ab88e3, 32'h42b3326b, 32'hc15af933, 32'hc281d729, 32'hc1f7122f};
test_label[1907] = '{32'hc15af933};
test_output[1907] = '{32'h42ce9193};
/*############ DEBUG ############
test_input[15256:15263] = '{18.3298529558, -35.2217124679, 77.5056331523, -85.7673572087, 89.5984763549, -13.6858392319, -64.920233262, -30.8838795546};
test_label[1907] = '{-13.6858392319};
test_output[1907] = '{103.284321186};
############ END DEBUG ############*/
test_input[15264:15271] = '{32'h425c669d, 32'h423a46a1, 32'hc27928e7, 32'hc2b3b31b, 32'hc1e37f33, 32'hc217d440, 32'hc1f9ac5b, 32'hc2161da9};
test_label[1908] = '{32'hc2b3b31b};
test_output[1908] = '{32'h4310f342};
/*############ DEBUG ############
test_input[15264:15271] = '{55.1002087009, 46.5689735529, -62.2899426389, -89.8498174306, -28.4371090912, -37.9572741375, -31.2091584614, -37.5289662746};
test_label[1908] = '{-89.8498174306};
test_output[1908] = '{144.950223323};
############ END DEBUG ############*/
test_input[15272:15279] = '{32'hc2bb8a65, 32'h407dc4ea, 32'h42497449, 32'hc1c80abf, 32'h41fe6c81, 32'h42990e2a, 32'h42b25cb0, 32'h424f3508};
test_label[1909] = '{32'h42b25cb0};
test_output[1909] = '{32'h3656882c};
/*############ DEBUG ############
test_input[15272:15279] = '{-93.7703048903, 3.96514356509, 50.3635591578, -25.0052476398, 31.8029802674, 76.5276650938, 89.1810316503, 51.8017890253};
test_label[1909] = '{89.1810316503};
test_output[1909] = '{3.19677472492e-06};
############ END DEBUG ############*/
test_input[15280:15287] = '{32'hc27e5b65, 32'h42561154, 32'h42ba1f11, 32'h4162da75, 32'h42a2ff57, 32'hc1bbc541, 32'h42a99965, 32'h41d1d028};
test_label[1910] = '{32'hc27e5b65};
test_output[1910] = '{32'h431ca673};
/*############ DEBUG ############
test_input[15280:15287] = '{-63.5892532471, 53.5169228453, 93.0606765386, 14.178334084, 81.4987099634, -23.4713158108, 84.7995958713, 26.2266383872};
test_label[1910] = '{-63.5892532471};
test_output[1910] = '{156.650197651};
############ END DEBUG ############*/
test_input[15288:15295] = '{32'hc207ffdc, 32'hbec48708, 32'h42c33f58, 32'h421d0711, 32'h42aad4ba, 32'h412ed248, 32'h410f611c, 32'h419b6c64};
test_label[1911] = '{32'h42c33f58};
test_output[1911] = '{32'h36a768a3};
/*############ DEBUG ############
test_input[15288:15295] = '{-33.9998609509, -0.383842715882, 97.6237167924, 39.25690139, 85.4154780877, 10.9263377318, 8.96120877238, 19.427925393};
test_label[1911] = '{97.6237167924};
test_output[1911] = '{4.98916897912e-06};
############ END DEBUG ############*/
test_input[15296:15303] = '{32'h42321316, 32'h4227e95b, 32'hc2c078d7, 32'hc28ac6cd, 32'hc2bc92e5, 32'h41ef5b7f, 32'hc2a4565f, 32'h425d076e};
test_label[1912] = '{32'h425d076e};
test_output[1912] = '{32'h37c44b3f};
/*############ DEBUG ############
test_input[15296:15303] = '{44.5186387291, 41.9778877523, -96.2360141712, -69.3882800616, -94.2869019365, 29.9196762184, -82.1686964638, 55.2572554364};
test_label[1912] = '{55.2572554364};
test_output[1912] = '{2.34000592856e-05};
############ END DEBUG ############*/
test_input[15304:15311] = '{32'h42189d7b, 32'hc278da09, 32'h429520c6, 32'hc109828e, 32'h428c7fea, 32'hc2a578c8, 32'h429617b3, 32'hc20c1faa};
test_label[1913] = '{32'h429520c6};
test_output[1913] = '{32'h3f77da77};
/*############ DEBUG ############
test_input[15304:15311] = '{38.1537909738, -62.2129260224, 74.5640096983, -8.59437398688, 70.2498351196, -82.7359023923, 75.0462894889, -35.0309231104};
test_label[1913] = '{74.5640096983};
test_output[1913] = '{0.968177241558};
############ END DEBUG ############*/
test_input[15312:15319] = '{32'h4064a3ab, 32'hc0bef9dd, 32'hc2bfc811, 32'hc23cd964, 32'h422661ae, 32'hc1a98a51, 32'h41232fa8, 32'hc2ad3ee0};
test_label[1914] = '{32'hc1a98a51};
test_output[1914] = '{32'h427b26d6};
/*############ DEBUG ############
test_input[15312:15319] = '{3.57248947731, -5.96800083252, -95.8907510072, -47.2122944371, 41.5953899629, -21.1925364018, 10.1991348671, -86.6228062516};
test_label[1914] = '{-21.1925364018};
test_output[1914] = '{62.7879263647};
############ END DEBUG ############*/
test_input[15320:15327] = '{32'hc298dac2, 32'h425c9a69, 32'h420f1804, 32'h413a1445, 32'hc20c3f24, 32'hc2b1aa98, 32'h4189b337, 32'hc22c46b9};
test_label[1915] = '{32'h413a1445};
test_output[1915] = '{32'h422e1558};
/*############ DEBUG ############
test_input[15320:15327] = '{-76.427259052, 55.1507916771, 35.7734514902, 11.6299486324, -35.0616616952, -88.8331879144, 17.2125066636, -43.069066436};
test_label[1915] = '{11.6299486324};
test_output[1915] = '{43.5208430485};
############ END DEBUG ############*/
test_input[15328:15335] = '{32'hc28283be, 32'h42bd5632, 32'h419dd9a8, 32'h40da3203, 32'h42595919, 32'h4266d08d, 32'hc0e63f1f, 32'hc2b94bb8};
test_label[1916] = '{32'h40da3203};
test_output[1916] = '{32'h42afb312};
/*############ DEBUG ############
test_input[15328:15335] = '{-65.2573104414, 94.6683521215, 19.7312767698, 6.8186050103, 54.3370090098, 57.7036616001, -7.1952050544, -92.64789102};
test_label[1916] = '{6.8186050103};
test_output[1916] = '{87.8497471112};
############ END DEBUG ############*/
test_input[15336:15343] = '{32'hc0b85f9d, 32'h42c57763, 32'hc201cb7c, 32'hc289658a, 32'hc20290e8, 32'h4281a1cd, 32'h411a93a7, 32'h41220fc6};
test_label[1917] = '{32'hc0b85f9d};
test_output[1917] = '{32'h42d0fd5d};
/*############ DEBUG ############
test_input[15336:15343] = '{-5.76167148802, 98.7331759007, -32.4487162346, -68.6983181177, -32.6415098886, 64.8160191167, 9.66104824183, 10.1288509987};
test_label[1917] = '{-5.76167148802};
test_output[1917] = '{104.494847389};
############ END DEBUG ############*/
test_input[15344:15351] = '{32'h4282a494, 32'hc2bd8bc2, 32'hc280ca19, 32'hc1ef38b2, 32'hc216df2d, 32'h419d694f, 32'hbf107ff4, 32'h42933856};
test_label[1918] = '{32'hc1ef38b2};
test_output[1918] = '{32'h42cf06a3};
/*############ DEBUG ############
test_input[15344:15351] = '{65.3214380816, -94.7729678272, -64.3947249556, -29.9026836149, -37.7179441612, 19.6764197328, -0.564452380822, 73.6100306516};
test_label[1918] = '{-29.9026836149};
test_output[1918] = '{103.512965603};
############ END DEBUG ############*/
test_input[15352:15359] = '{32'hc09785ec, 32'hc214ea5a, 32'hc29f6cef, 32'hc22e5c94, 32'h426539b3, 32'h3ef264dc, 32'h42700e1d, 32'hc2a9cb5e};
test_label[1919] = '{32'h426539b3};
test_output[1919] = '{32'h403168a6};
/*############ DEBUG ############
test_input[15352:15359] = '{-4.73509791159, -37.2288597689, -79.7127571488, -43.5904075897, 57.3063478158, 0.473425734797, 60.0137830379, -84.8972030637};
test_label[1919] = '{57.3063478158};
test_output[1919] = '{2.7720121905};
############ END DEBUG ############*/
test_input[15360:15367] = '{32'h42bc9533, 32'h424250bb, 32'hc288285b, 32'h4201d93a, 32'h4154095d, 32'h4291c2cc, 32'h420ac0a6, 32'hc1e97c93};
test_label[1920] = '{32'h42bc9533};
test_output[1920] = '{32'h300a3168};
/*############ DEBUG ############
test_input[15360:15367] = '{94.2914019973, 48.5788388971, -68.0788198036, 32.4621338322, 13.2522862911, 72.8804601929, 34.6881331964, -29.1858272124};
test_label[1920] = '{94.2914019973};
test_output[1920] = '{5.02743180546e-10};
############ END DEBUG ############*/
test_input[15368:15375] = '{32'h429aa506, 32'hc217848e, 32'h42483d22, 32'hbf8d9b43, 32'hc2a5841d, 32'h424779e7, 32'h4296121b, 32'hc203030e};
test_label[1921] = '{32'h424779e7};
test_output[1921] = '{32'h41dc666a};
/*############ DEBUG ############
test_input[15368:15375] = '{77.3223106636, -37.8794487837, 50.0597015365, -1.1063006679, -82.7580368558, 49.8690463257, 75.0353595503, -32.7529842351};
test_label[1921] = '{49.8690463257};
test_output[1921] = '{27.5500059318};
############ END DEBUG ############*/
test_input[15376:15383] = '{32'h429ded0c, 32'h42ba6fae, 32'hc1dc7c24, 32'h4240399c, 32'h42a93e7f, 32'hc14b2b70, 32'hc2939e47, 32'h42a602ea};
test_label[1922] = '{32'hc2939e47};
test_output[1922] = '{32'h43270709};
/*############ DEBUG ############
test_input[15376:15383] = '{78.9629829716, 93.2181244045, -27.5606147846, 48.0562598056, 84.6220652281, -12.6981050491, -73.8091317784, 83.0056920393};
test_label[1922] = '{-73.8091317784};
test_output[1922] = '{167.027478346};
############ END DEBUG ############*/
test_input[15384:15391] = '{32'hc27a7a54, 32'hc293f8ea, 32'hc2aa595a, 32'hc2c548f3, 32'hc24a6dd0, 32'h426cb564, 32'h42780e6d, 32'h42a8b3a9};
test_label[1923] = '{32'hc27a7a54};
test_output[1923] = '{32'h4312f86a};
/*############ DEBUG ############
test_input[15384:15391] = '{-62.6194625544, -73.9861619258, -85.1745163717, -98.642479569, -50.6072406769, 59.1771386255, 62.0140877993, 84.3509013664};
test_label[1923] = '{-62.6194625544};
test_output[1923] = '{146.970363921};
############ END DEBUG ############*/
test_input[15392:15399] = '{32'hc0ce82ab, 32'h4295b8c4, 32'h40c905ea, 32'hc28d8ae6, 32'h40d3cb9b, 32'hc1f1390a, 32'hc18e2fc2, 32'hc11f6aee};
test_label[1924] = '{32'hc11f6aee};
test_output[1924] = '{32'h42a9a622};
/*############ DEBUG ############
test_input[15392:15399] = '{-6.45345064564, 74.8608717481, 6.28197199602, -70.7712867409, 6.61860409623, -30.1528515837, -17.7733188992, -9.96360567321};
test_label[1924] = '{-9.96360567321};
test_output[1924] = '{84.8244774213};
############ END DEBUG ############*/
test_input[15400:15407] = '{32'hc21e6b61, 32'hc1eb391a, 32'hc22ded78, 32'h41e28898, 32'hc005e6e2, 32'hbd55727d, 32'h428b4634, 32'h405e5db4};
test_label[1925] = '{32'hc21e6b61};
test_output[1925] = '{32'h42da7be4};
/*############ DEBUG ############
test_input[15400:15407] = '{-39.6048604195, -29.4028818517, -43.481904055, 28.3166965793, -2.0922169334, -0.0521111378686, 69.6371164493, 3.47446913307};
test_label[1925] = '{-39.6048604195};
test_output[1925] = '{109.241976869};
############ END DEBUG ############*/
test_input[15408:15415] = '{32'h41c838f0, 32'hc04a97b8, 32'hc2a0116c, 32'hc2c66704, 32'hc29db1b0, 32'h4085545b, 32'hc2af62fc, 32'h429f0b90};
test_label[1926] = '{32'hc04a97b8};
test_output[1926] = '{32'h42a5604d};
/*############ DEBUG ############
test_input[15408:15415] = '{25.0278011575, -3.16551007364, -80.0340305004, -99.2012007528, -78.8470487681, 4.1665472921, -87.6933278577, 79.5225797651};
test_label[1926] = '{-3.16551007364};
test_output[1926] = '{82.6880898387};
############ END DEBUG ############*/
test_input[15416:15423] = '{32'h425590f5, 32'hc2b45522, 32'hc262a6da, 32'h3fa6c0b0, 32'hc256e336, 32'h417a8f9e, 32'hc290c05c, 32'hc2a215dd};
test_label[1927] = '{32'h425590f5};
test_output[1927] = '{32'h80000000};
/*############ DEBUG ############
test_input[15416:15423] = '{53.3915588774, -90.1662722022, -56.662942809, 1.30275539732, -53.7218874474, 15.6600630603, -72.3757042837, -81.0427049028};
test_label[1927] = '{53.3915588774};
test_output[1927] = '{-0.0};
############ END DEBUG ############*/
test_input[15424:15431] = '{32'h42094615, 32'h415a2b58, 32'hc2b4e687, 32'h42c773d1, 32'hc20b7c0e, 32'hc023eda2, 32'hc224983d, 32'hc12c788e};
test_label[1928] = '{32'hc023eda2};
test_output[1928] = '{32'h42cc933e};
/*############ DEBUG ############
test_input[15424:15431] = '{34.318439991, 13.6355822278, -90.4502484468, 99.7262023972, -34.8711462317, -2.56137892703, -41.1486720906, -10.7794325811};
test_label[1928] = '{-2.56137892703};
test_output[1928] = '{102.287581324};
############ END DEBUG ############*/
test_input[15432:15439] = '{32'hc25fdd3c, 32'hc22ac946, 32'h41873e66, 32'hc211fa01, 32'hc26c70fc, 32'hc2a55133, 32'hc27a92bd, 32'h42b792e3};
test_label[1929] = '{32'hc2a55133};
test_output[1929] = '{32'h432e720b};
/*############ DEBUG ############
test_input[15432:15439] = '{-55.9660495054, -42.6965551454, 16.9054673132, -36.4941429181, -59.1103358093, -82.6585941927, -62.6433001004, 91.7868910273};
test_label[1929] = '{-82.6585941927};
test_output[1929] = '{174.44548522};
############ END DEBUG ############*/
test_input[15440:15447] = '{32'h426183f5, 32'h40064f6c, 32'hc191fb25, 32'h4114bbec, 32'hc20b597d, 32'hc2941693, 32'hc1ced22b, 32'hc28ab8e9};
test_label[1930] = '{32'hc2941693};
test_output[1930] = '{32'h43026c47};
/*############ DEBUG ############
test_input[15440:15447] = '{56.378864858, 2.09859757624, -18.2476294956, 9.29587924417, -34.8373916606, -74.0440905335, -25.8526211835, -69.3611522847};
test_label[1930] = '{-74.0440905335};
test_output[1930] = '{130.422955392};
############ END DEBUG ############*/
test_input[15448:15455] = '{32'hc1512fd8, 32'hc14e1fea, 32'hc29ac4a1, 32'hc1398b2f, 32'h42a7f063, 32'h4038c8c7, 32'h42b1bb36, 32'h42c39475};
test_label[1931] = '{32'hc1398b2f};
test_output[1931] = '{32'h42dac5ec};
/*############ DEBUG ############
test_input[15448:15455] = '{-13.0741804019, -12.8827914957, -77.3840372227, -11.5964802176, 83.9695076876, 2.88725437177, 88.8656436851, 97.7899526946};
test_label[1931] = '{-11.5964802176};
test_output[1931] = '{109.386567012};
############ END DEBUG ############*/
test_input[15456:15463] = '{32'hc1a65156, 32'h41da7099, 32'h419d3db1, 32'hc2a4dd1e, 32'h4258b2ea, 32'h426a6a03, 32'hc2c08b94, 32'h426f2543};
test_label[1932] = '{32'h4258b2ea};
test_output[1932] = '{32'h40bc372f};
/*############ DEBUG ############
test_input[15456:15463] = '{-20.7897143854, 27.3049791967, 19.6551220381, -82.4318692586, 54.1747208417, 58.6035282122, -96.2726116013, 59.7863866706};
test_label[1932] = '{54.1747208417};
test_output[1932] = '{5.8817361904};
############ END DEBUG ############*/
test_input[15464:15471] = '{32'h424f8a69, 32'h42bb18d0, 32'h42a470c0, 32'hc258d83a, 32'hc1e5cda1, 32'h42848a3f, 32'h42bbae50, 32'h4158da01};
test_label[1933] = '{32'h424f8a69};
test_output[1933] = '{32'h422a0d61};
/*############ DEBUG ############
test_input[15464:15471] = '{51.8851679166, 93.5484647622, 82.2202143805, -54.2111606505, -28.7254052994, 66.2700120035, 93.8404562873, 13.5532239282};
test_label[1933] = '{51.8851679166};
test_output[1933] = '{42.5130646662};
############ END DEBUG ############*/
test_input[15472:15479] = '{32'hc24996d8, 32'h42a4a293, 32'hc29e325b, 32'hc2bde440, 32'hc18555f8, 32'hc16ef415, 32'hc230d0cd, 32'h418c0277};
test_label[1934] = '{32'h418c0277};
test_output[1934] = '{32'h4281a1f5};
/*############ DEBUG ############
test_input[15472:15479] = '{-50.3973085235, 82.3175247362, -79.0983529761, -94.9457993056, -16.6669761069, -14.9345904426, -44.2039068125, 17.5012031204};
test_label[1934] = '{17.5012031204};
test_output[1934] = '{64.8163216158};
############ END DEBUG ############*/
test_input[15480:15487] = '{32'h429fc711, 32'h4295d326, 32'h429ecf27, 32'hc282901f, 32'hbeab4da6, 32'hc121b7e5, 32'hc2580ac2, 32'h42c2c9dc};
test_label[1935] = '{32'hc2580ac2};
test_output[1935] = '{32'h4317679e};
/*############ DEBUG ############
test_input[15480:15487] = '{79.8888053509, 74.9124014727, 79.4045917661, -65.2814845523, -0.334576797623, -10.107396406, -54.0105042286, 97.3942545509};
test_label[1935] = '{-54.0105042286};
test_output[1935] = '{151.40475882};
############ END DEBUG ############*/
test_input[15488:15495] = '{32'hc29a68f6, 32'h3d0c358f, 32'h422a607b, 32'hc232055a, 32'hc1d57670, 32'h41881672, 32'hc2a8dbb1, 32'hc2c795f1};
test_label[1936] = '{32'hc2c795f1};
test_output[1936] = '{32'h430e6317};
/*############ DEBUG ############
test_input[15488:15495] = '{-77.2049996684, 0.0342307631226, 42.5942202688, -44.5052274763, -26.6828312843, 17.010959859, -84.4290857596, -99.792856175};
test_label[1936] = '{-99.792856175};
test_output[1936] = '{142.387076444};
############ END DEBUG ############*/
test_input[15496:15503] = '{32'h42b83d6e, 32'h42772266, 32'h4234692b, 32'h42a5ee31, 32'h41e476a4, 32'hc0bf95a2, 32'hc2ba75f6, 32'h41ad3a06};
test_label[1937] = '{32'h42b83d6e};
test_output[1937] = '{32'h38ddb031};
/*############ DEBUG ############
test_input[15496:15503] = '{92.1199806015, 61.7835913459, 45.1027012597, 82.9652147772, 28.5579303087, -5.98701561553, -93.2303926494, 21.6533318779};
test_label[1937] = '{92.1199806015};
test_output[1937] = '{0.000105709194859};
############ END DEBUG ############*/
test_input[15504:15511] = '{32'hc2aaa6b3, 32'h41599ff3, 32'hc259f5e6, 32'hc1d75991, 32'h410e2426, 32'h42b9d3dc, 32'h41ac5990, 32'h42916c34};
test_label[1938] = '{32'h42b9d3dc};
test_output[1938] = '{32'h30e75d62};
/*############ DEBUG ############
test_input[15504:15511] = '{-85.325581843, 13.6015500452, -54.4901348546, -26.9187341329, 8.88382498521, 92.9137842759, 21.5437317013, 72.7113341805};
test_label[1938] = '{92.9137842759};
test_output[1938] = '{1.68340030946e-09};
############ END DEBUG ############*/
test_input[15512:15519] = '{32'hc0fed85a, 32'hc2a08a25, 32'hc23c076c, 32'h41c02d04, 32'hc22f46e3, 32'h4226113c, 32'hc2a54f12, 32'hc16de4fc};
test_label[1939] = '{32'hc2a08a25};
test_output[1939] = '{32'h42f392c3};
/*############ DEBUG ############
test_input[15512:15519] = '{-7.96391007862, -80.2698123546, -47.0072461943, 24.0219807987, -43.8192242907, 41.5168293342, -82.6544363952, -14.8684039252};
test_label[1939] = '{-80.2698123546};
test_output[1939] = '{121.786641714};
############ END DEBUG ############*/
test_input[15520:15527] = '{32'hc182c755, 32'h424372c6, 32'hc237cf02, 32'h4248ca5d, 32'hc2415a0b, 32'hc0c17fa7, 32'h42b2dec1, 32'hc25e9f33};
test_label[1940] = '{32'h4248ca5d};
test_output[1940] = '{32'h421cf325};
/*############ DEBUG ############
test_input[15520:15527] = '{-16.347330963, 48.8620851831, -45.9521549598, 50.1976217901, -48.3379313104, -6.04683241505, 89.435067291, -55.6554679721};
test_label[1940] = '{50.1976217901};
test_output[1940] = '{39.2374455009};
############ END DEBUG ############*/
test_input[15528:15535] = '{32'hc262164e, 32'h41a87da6, 32'hc2bd1321, 32'h4288ea0c, 32'h42731f9e, 32'hc181f64c, 32'h41859057, 32'hc23abf44};
test_label[1941] = '{32'hc23abf44};
test_output[1941] = '{32'h42e649eb};
/*############ DEBUG ############
test_input[15528:15535] = '{-56.5217830083, 21.0613509146, -94.5373641589, 68.4571261947, 60.7808752809, -16.245261887, 16.6954787787, -46.6867811017};
test_label[1941] = '{-46.6867811017};
test_output[1941] = '{115.144370899};
############ END DEBUG ############*/
test_input[15536:15543] = '{32'hc1d3ad36, 32'hc0ff8c3a, 32'hc147f8ad, 32'h4098c640, 32'hc28876d3, 32'hc19f1012, 32'h41c10734, 32'h420bb6cd};
test_label[1942] = '{32'hc19f1012};
test_output[1942] = '{32'h425b3edc};
/*############ DEBUG ############
test_input[15536:15543] = '{-26.4595748167, -7.98586750439, -12.498212055, 4.77420061008, -68.2320756931, -19.8828471034, 24.1285164199, 34.9285173443};
test_label[1942] = '{-19.8828471034};
test_output[1942] = '{54.8113848469};
############ END DEBUG ############*/
test_input[15544:15551] = '{32'h42807bb7, 32'hc2396f58, 32'hc2348dec, 32'hc2821417, 32'hc1312968, 32'h428d5677, 32'h41d5dea8, 32'hc2388b82};
test_label[1943] = '{32'h41d5dea8};
test_output[1943] = '{32'h422fbf41};
/*############ DEBUG ############
test_input[15544:15551] = '{64.241627286, -46.3587323991, -45.1385957242, -65.0392416249, -11.0726088295, 70.668873076, 26.733718891, -46.1362363755};
test_label[1943] = '{26.733718891};
test_output[1943] = '{43.9367697773};
############ END DEBUG ############*/
test_input[15552:15559] = '{32'h429b695d, 32'hc18bb4d8, 32'hc0133008, 32'h42a7a71b, 32'h42c2f98c, 32'h41c4bb13, 32'h422fd436, 32'hc1b72c90};
test_label[1944] = '{32'hc18bb4d8};
test_output[1944] = '{32'h42e5e6c2};
/*############ DEBUG ############
test_input[15552:15559] = '{77.7057842335, -17.4633033013, -2.29980659339, 83.8263787747, 97.4873950925, 24.5913445254, 43.9572386998, -22.8967583878};
test_label[1944] = '{-17.4633033013};
test_output[1944] = '{114.950699563};
############ END DEBUG ############*/
test_input[15560:15567] = '{32'hc12c2d47, 32'h4018fa93, 32'hc260a782, 32'h42ae9570, 32'hc28518f2, 32'h42b07371, 32'hc0c7c9af, 32'h41012c87};
test_label[1945] = '{32'hc0c7c9af};
test_output[1945] = '{32'h42bd99cd};
/*############ DEBUG ############
test_input[15560:15567] = '{-10.7610539729, 2.39029372076, -56.163581186, 87.2918664272, -66.5487187762, 88.2254679527, -6.24336965587, 8.07337126403};
test_label[1945] = '{-6.24336965587};
test_output[1945] = '{94.8003944063};
############ END DEBUG ############*/
test_input[15568:15575] = '{32'h41c749cf, 32'hc0810f30, 32'h4275cc0d, 32'h42aaab33, 32'h42a00376, 32'hc285d45a, 32'h418b2d00, 32'hc2b6e984};
test_label[1946] = '{32'h42aaab33};
test_output[1946] = '{32'h3b9eb9ae};
/*############ DEBUG ############
test_input[15568:15575] = '{24.9110396081, -4.03310392567, 61.4492676633, 85.3343709946, 80.0067613432, -66.9147489318, 17.396973248, -91.4560868631};
test_label[1946] = '{85.3343709946};
test_output[1946] = '{0.0048439122122};
############ END DEBUG ############*/
test_input[15576:15583] = '{32'h4213b3f0, 32'h427862e6, 32'h3f1bde0b, 32'h41c0576d, 32'h428f1c6a, 32'hc1b865d2, 32'hc19476c6, 32'hc134e1dd};
test_label[1947] = '{32'hc19476c6};
test_output[1947] = '{32'h42b43a26};
/*############ DEBUG ############
test_input[15576:15583] = '{36.9257198125, 62.0965817985, 0.608856840934, 24.0426885495, 71.5554963193, -23.0497162431, -18.5579940365, -11.305142359};
test_label[1947] = '{-18.5579940365};
test_output[1947] = '{90.113568344};
############ END DEBUG ############*/
test_input[15584:15591] = '{32'hc2bf33c2, 32'h41a47754, 32'hc0d08cdb, 32'hc205f8a2, 32'hc284d20e, 32'hc25a17e0, 32'h421f4a18, 32'hc1d82f6a};
test_label[1948] = '{32'hc0d08cdb};
test_output[1948] = '{32'h42395bb3};
/*############ DEBUG ############
test_input[15584:15591] = '{-95.6010927508, 20.5582665924, -6.51719423263, -33.4928065171, -66.410265295, -54.5233157633, 39.8223572022, -27.0231506295};
test_label[1948] = '{-6.51719423263};
test_output[1948] = '{46.3395514391};
############ END DEBUG ############*/
test_input[15592:15599] = '{32'hc263281a, 32'hc2ad857a, 32'h429b91eb, 32'hc2001814, 32'hc2bbf1e0, 32'hc178df3f, 32'h42910a8b, 32'h40a0ce6d};
test_label[1949] = '{32'hc263281a};
test_output[1949] = '{32'h4306944e};
/*############ DEBUG ############
test_input[15592:15599] = '{-56.7891610944, -86.7606951565, 77.7849981125, -32.023513958, -93.9724133021, -15.5545030747, 72.5205882425, 5.02519833546};
test_label[1949] = '{-56.7891610944};
test_output[1949] = '{134.57931832};
############ END DEBUG ############*/
test_input[15600:15607] = '{32'hc252cc1f, 32'h41d66fca, 32'hc2b64488, 32'h429e19b5, 32'hc297b43b, 32'hc2c60395, 32'h428ef37f, 32'h41f2839c};
test_label[1950] = '{32'h41f2839c};
test_output[1950] = '{32'h4242f223};
/*############ DEBUG ############
test_input[15600:15607] = '{-52.6993374298, 26.8045853135, -91.1338502809, 79.0502089522, -75.8520119136, -99.0069984139, 71.4755808131, 30.3142618798};
test_label[1950] = '{30.3142618798};
test_output[1950] = '{48.736460252};
############ END DEBUG ############*/
test_input[15608:15615] = '{32'hc031c616, 32'hc119a031, 32'h42962c27, 32'h428d81da, 32'h42c1a98a, 32'h42aa8d82, 32'hc2329d19, 32'h41bbc7e5};
test_label[1951] = '{32'h42aa8d82};
test_output[1951] = '{32'h4138e049};
/*############ DEBUG ############
test_input[15608:15615] = '{-2.7777151804, -9.60160955876, 75.0862373329, 70.753617922, 96.8311316201, 85.276383623, -44.6534174272, 23.4726041301};
test_label[1951] = '{85.276383623};
test_output[1951] = '{11.5547575879};
############ END DEBUG ############*/
test_input[15616:15623] = '{32'hc227b0e4, 32'hc2a0ee0a, 32'hc273c90d, 32'hc02e88db, 32'hc2492d3f, 32'h42a08352, 32'h41acc9bc, 32'hc299fdee};
test_label[1952] = '{32'hc2492d3f};
test_output[1952] = '{32'h43028cf9};
/*############ DEBUG ############
test_input[15616:15623] = '{-41.9227454201, -80.4649171974, -60.9463402414, -2.7271030948, -50.2941864965, 80.2564834386, 21.5985038438, -76.9959593865};
test_label[1952] = '{-50.2941864965};
test_output[1952] = '{130.550669935};
############ END DEBUG ############*/
test_input[15624:15631] = '{32'hc2ad1bdc, 32'hc282a5ac, 32'hc29ec197, 32'hc2ab6b0c, 32'h41cd0299, 32'hc24a44b4, 32'h42736786, 32'hc1f4f823};
test_label[1953] = '{32'h42736786};
test_output[1953] = '{32'h26200000};
/*############ DEBUG ############
test_input[15624:15631] = '{-86.5544118433, -65.3235771132, -79.378107363, -85.7090765258, 25.6262687345, -50.567091502, 60.8510964909, -30.6211611391};
test_label[1953] = '{60.8510964909};
test_output[1953] = '{5.55111512313e-16};
############ END DEBUG ############*/
test_input[15632:15639] = '{32'h42837abb, 32'h3e06b358, 32'h421fc7e3, 32'h4159deab, 32'hc27d424d, 32'hc0e9097d, 32'h4293c0c2, 32'h41fbc6a2};
test_label[1954] = '{32'hc27d424d};
test_output[1954] = '{32'h43093107};
/*############ DEBUG ############
test_input[15632:15639] = '{65.739709682, 0.131543516918, 39.9452019793, 13.6168626412, -63.3147483822, -7.282408039, 73.8764765757, 31.4719893217};
test_label[1954] = '{-63.3147483822};
test_output[1954] = '{137.191517497};
############ END DEBUG ############*/
test_input[15640:15647] = '{32'h4288fb45, 32'hc2252b8e, 32'hc1ff7d6f, 32'h4251fdac, 32'hc2478fc2, 32'h41fa04e7, 32'h418bb96c, 32'h42b8a324};
test_label[1955] = '{32'hc1ff7d6f};
test_output[1955] = '{32'h42f88280};
/*############ DEBUG ############
test_input[15640:15647] = '{68.4907636686, -41.2925351356, -31.9362470726, 52.4977259912, -49.8903870646, 31.252393097, 17.465538164, 92.318637193};
test_label[1955] = '{-31.9362470726};
test_output[1955] = '{124.254884266};
############ END DEBUG ############*/
test_input[15648:15655] = '{32'hc28680f5, 32'h41e4f004, 32'hc264b749, 32'h42bbaf1a, 32'hc2a72479, 32'hc23f4d27, 32'hc2609024, 32'h42102e1a};
test_label[1956] = '{32'hc23f4d27};
test_output[1956] = '{32'h430daad7};
/*############ DEBUG ############
test_input[15648:15655] = '{-67.2518698717, 28.6171952132, -57.1789887691, 93.8419948989, -83.5712362717, -47.8253453966, -56.1407615233, 36.0450218501};
test_label[1956] = '{-47.8253453966};
test_output[1956] = '{141.667340296};
############ END DEBUG ############*/
test_input[15656:15663] = '{32'h4209b9ca, 32'hc16792f2, 32'hc289f1f3, 32'hc2448b8d, 32'h42898673, 32'h4280d614, 32'h42bd46d4, 32'h4262ee7e};
test_label[1957] = '{32'h42bd46d4};
test_output[1957] = '{32'h2cce3000};
/*############ DEBUG ############
test_input[15656:15663] = '{34.4314332691, -14.4733754868, -68.9725580848, -49.1362811575, 68.7625969359, 64.4181217682, 94.6383392633, 56.732901245};
test_label[1957] = '{94.6383392633};
test_output[1957] = '{5.8602012132e-12};
############ END DEBUG ############*/
test_input[15664:15671] = '{32'h42533c97, 32'h40e53f01, 32'h427f76b1, 32'hc279fd87, 32'h42af4047, 32'hc0e1f6b4, 32'h41c4b37a, 32'h423ec3a3};
test_label[1958] = '{32'h42af4047};
test_output[1958] = '{32'h2e532640};
/*############ DEBUG ############
test_input[15664:15671] = '{52.8091711699, 7.16394098945, 63.8659091891, -62.4975846724, 87.6255394075, -7.06136510537, 24.587635174, 47.6910501617};
test_label[1958] = '{87.6255394075};
test_output[1958] = '{4.80098183442e-11};
############ END DEBUG ############*/
test_input[15672:15679] = '{32'hc2949e4d, 32'hc11117bf, 32'h3f378d7e, 32'hc1f90a65, 32'h425910be, 32'hc27d0d89, 32'h3fd18533, 32'hc1ca7b2f};
test_label[1959] = '{32'hc11117bf};
test_output[1959] = '{32'h427d56ae};
/*############ DEBUG ############
test_input[15672:15679] = '{-74.3091820433, -9.0682976058, 0.717002756769, -31.1300749741, 54.2663499157, -63.2632177536, 1.63687747618, -25.3101481885};
test_label[1959] = '{-9.0682976058};
test_output[1959] = '{63.3346475215};
############ END DEBUG ############*/
test_input[15680:15687] = '{32'hc1c45603, 32'h41e8780d, 32'hc2667f4e, 32'h42a68d27, 32'hc261263b, 32'h426de58f, 32'h42167672, 32'hc2c1c7a7};
test_label[1960] = '{32'h42a68d27};
test_output[1960] = '{32'h2e4a7ca0};
/*############ DEBUG ############
test_input[15680:15687] = '{-24.5419983952, 29.0586178153, -57.6243221445, 83.2756867237, -56.2873338611, 59.4741782987, 37.6156707936, -96.8899486405};
test_label[1960] = '{83.2756867237};
test_output[1960] = '{4.60401716761e-11};
############ END DEBUG ############*/
test_input[15688:15695] = '{32'hc1d21a26, 32'hc2a9ec1d, 32'hc23aea07, 32'hc170d357, 32'hc216d4b2, 32'hc19bf6a6, 32'hc1fbdbb7, 32'h42888442};
test_label[1961] = '{32'hc1fbdbb7};
test_output[1961] = '{32'h42c77b30};
/*############ DEBUG ############
test_input[15688:15695] = '{-26.2627683068, -84.9611610089, -46.7285405435, -15.0515969969, -37.7077112119, -19.4954339847, -31.4822818361, 68.2583171303};
test_label[1961] = '{-31.4822818361};
test_output[1961] = '{99.7405989663};
############ END DEBUG ############*/
test_input[15696:15703] = '{32'hc2139be9, 32'hc202980e, 32'h405afcdc, 32'hbead8b75, 32'h42a2381d, 32'h42a492e1, 32'hc28df983, 32'h42af0709};
test_label[1962] = '{32'hc28df983};
test_output[1962] = '{32'h431e8211};
/*############ DEBUG ############
test_input[15696:15703] = '{-36.9022561308, -32.6484921599, 3.42168339768, -0.338954609605, 81.1095949904, 82.286874174, -70.9873282517, 87.513740792};
test_label[1962] = '{-70.9873282517};
test_output[1962] = '{158.508069493};
############ END DEBUG ############*/
test_input[15704:15711] = '{32'h42296bf9, 32'hc29eafca, 32'h42738eec, 32'hc287f38f, 32'h42a8ef62, 32'h425c1f50, 32'h4198bc64, 32'h42a82a72};
test_label[1963] = '{32'h42a82a72};
test_output[1963] = '{32'h3f67628b};
/*############ DEBUG ############
test_input[15704:15711] = '{42.3554404691, -79.3433369046, 60.8895720826, -67.9757007227, 84.4675430896, 55.030579514, 19.0919870064, 84.082903729};
test_label[1963] = '{84.082903729};
test_output[1963] = '{0.90384740025};
############ END DEBUG ############*/
test_input[15712:15719] = '{32'hc2aa8ea5, 32'h41af5949, 32'h42aabda0, 32'hc237a049, 32'h42ad4bc6, 32'hc2a48e1d, 32'h4202dee1, 32'h421d1c86};
test_label[1964] = '{32'h421d1c86};
test_output[1964] = '{32'h423e76c5};
/*############ DEBUG ############
test_input[15712:15719] = '{-85.2786013881, 21.9185955277, 85.370363983, -45.9065275974, 86.6479973104, -82.2775688082, 32.7176543877, 39.2778538107};
test_label[1964] = '{39.2778538107};
test_output[1964] = '{47.6159843888};
############ END DEBUG ############*/
test_input[15720:15727] = '{32'hc202049f, 32'hc1fb574e, 32'hc212e201, 32'h428bf38e, 32'hc2076cf1, 32'hc2374623, 32'hc28c951e, 32'hc20c1219};
test_label[1965] = '{32'hc2076cf1};
test_output[1965] = '{32'h42cfaa07};
/*############ DEBUG ############
test_input[15720:15727] = '{-32.5045122362, -31.4176289066, -36.7207082154, 69.9756943009, -33.856387284, -45.8184917346, -70.2912473065, -35.0176736073};
test_label[1965] = '{-33.856387284};
test_output[1965] = '{103.832081585};
############ END DEBUG ############*/
test_input[15728:15735] = '{32'hc2b866b9, 32'h425cca70, 32'h429c2dd3, 32'hc21d5e0b, 32'hc29a08ab, 32'hc2ae7dc0, 32'hc2c52863, 32'h414b37e5};
test_label[1966] = '{32'h425cca70};
test_output[1966] = '{32'h41b7226a};
/*############ DEBUG ############
test_input[15728:15735] = '{-92.2006302105, 55.1976931603, 78.0894971582, -39.3418382573, -77.0169294044, -87.2456088972, -98.578878975, 12.7011457403};
test_label[1966] = '{55.1976931603};
test_output[1966] = '{22.891803998};
############ END DEBUG ############*/
test_input[15736:15743] = '{32'hc2b249cf, 32'hc187cfae, 32'h428a9dc4, 32'hc24f35f9, 32'hc24316f7, 32'hc13945a2, 32'h410b5ed7, 32'h429867f5};
test_label[1967] = '{32'hc24316f7};
test_output[1967] = '{32'h42f9f3f5};
/*############ DEBUG ############
test_input[15736:15743] = '{-89.1441558565, -16.9764053051, 69.3081376395, -51.8027083928, -48.7724273238, -11.5795005173, 8.71065446636, 76.2030404017};
test_label[1967] = '{-48.7724273238};
test_output[1967] = '{124.976480148};
############ END DEBUG ############*/
test_input[15744:15751] = '{32'hc2ac7ee8, 32'h42a67aa6, 32'hc1b09d31, 32'h425f2f84, 32'h425fe812, 32'h42526be2, 32'hc2172ec2, 32'hc270aba2};
test_label[1968] = '{32'hc2172ec2};
test_output[1968] = '{32'h42f21207};
/*############ DEBUG ############
test_input[15744:15751] = '{-86.2478620518, 83.2395483227, -22.0767532153, 55.7964030886, 55.9766321625, 52.6053545384, -37.795660954, -60.1676107802};
test_label[1968] = '{-37.795660954};
test_output[1968] = '{121.035209277};
############ END DEBUG ############*/
test_input[15752:15759] = '{32'hc2a6f22b, 32'h420476c2, 32'h428e53f2, 32'hc07878c2, 32'h422abd1f, 32'hc197d8e8, 32'h42736d9e, 32'hc297d262};
test_label[1969] = '{32'h422abd1f};
test_output[1969] = '{32'h41e3d59d};
/*############ DEBUG ############
test_input[15752:15759] = '{-83.4729858877, 33.1159732439, 71.163957097, -3.88237053767, 42.6846867425, -18.9809117841, 60.8570496172, -75.9109049253};
test_label[1969] = '{42.6846867425};
test_output[1969] = '{28.4793037556};
############ END DEBUG ############*/
test_input[15760:15767] = '{32'hc13c6009, 32'hc2920660, 32'h423cc5b4, 32'hc1559b53, 32'hc201de29, 32'h41ee3a56, 32'h42c38e07, 32'hc2c327d3};
test_label[1970] = '{32'h423cc5b4};
test_output[1970] = '{32'h424a565a};
/*############ DEBUG ############
test_input[15760:15767] = '{-11.7734460226, -73.0124525587, 47.1930704968, -13.3504210667, -32.4669533119, 29.7784842281, 97.777399997, -97.5777789874};
test_label[1970] = '{47.1930704968};
test_output[1970] = '{50.5843295002};
############ END DEBUG ############*/
test_input[15768:15775] = '{32'h4270a4ed, 32'h42ac2f1c, 32'hc2c756b3, 32'h4190d2db, 32'h42a295c8, 32'hc2287865, 32'h42a5edd8, 32'hc21bcdd8};
test_label[1971] = '{32'hc2287865};
test_output[1971] = '{32'h430042a5};
/*############ DEBUG ############
test_input[15768:15775] = '{60.1610613469, 86.0920106312, -99.6693336571, 18.1029572874, 81.2925405894, -42.1175710144, 82.9645418532, -38.9510209419};
test_label[1971] = '{-42.1175710144};
test_output[1971] = '{128.260334365};
############ END DEBUG ############*/
test_input[15776:15783] = '{32'h40c39d4b, 32'h42c4916c, 32'h42a14d8d, 32'h42352f1e, 32'h4214f90a, 32'h429eda6f, 32'hc1ec71a5, 32'hc22c97cb};
test_label[1972] = '{32'h42352f1e};
test_output[1972] = '{32'h4253f3ba};
/*############ DEBUG ############
test_input[15776:15783] = '{6.11295100652, 98.2840248167, 80.6514628497, 45.2960110096, 37.2432013218, 79.4266291351, -29.5554905981, -43.1482337044};
test_label[1972] = '{45.2960110096};
test_output[1972] = '{52.9880138355};
############ END DEBUG ############*/
test_input[15784:15791] = '{32'hc023b230, 32'hc129fe5c, 32'hc1338eec, 32'h4283e09c, 32'h42a0d8e2, 32'h40360743, 32'h429f4ed5, 32'hc27b3af9};
test_label[1973] = '{32'hc129fe5c};
test_output[1973] = '{32'h42b6db8e};
/*############ DEBUG ############
test_input[15784:15791] = '{-2.55775060074, -10.6245998631, -11.2223930945, 65.9386935632, 80.4236009024, 2.84419333869, 79.6539681601, -62.807591261};
test_label[1973] = '{-10.6245998631};
test_output[1973] = '{91.4288154139};
############ END DEBUG ############*/
test_input[15792:15799] = '{32'h42aa225a, 32'h4174f377, 32'h42099ffb, 32'hc26e1b36, 32'h409054d6, 32'h4187836b, 32'h426ab623, 32'hc184861e};
test_label[1974] = '{32'h42099ffb};
test_output[1974] = '{32'h424aa4ba};
/*############ DEBUG ############
test_input[15792:15799] = '{85.0670963797, 15.3094393207, 34.4062292641, -59.5265731629, 4.51035590647, 16.9391686168, 58.6778676861, -16.5654874481};
test_label[1974] = '{34.4062292641};
test_output[1974] = '{50.6608671156};
############ END DEBUG ############*/
test_input[15800:15807] = '{32'h42712ff8, 32'h42957c6f, 32'hc1972645, 32'h42b0806d, 32'h423a15a3, 32'h42a26113, 32'h42c523d4, 32'h42ab2644};
test_label[1975] = '{32'h42c523d4};
test_output[1975] = '{32'h381408ba};
/*############ DEBUG ############
test_input[15800:15807] = '{60.2968462035, 74.7430331301, -18.8936869854, 88.2508314948, 46.5211308623, 81.1896008937, 98.5699788203, 85.5747395961};
test_label[1975] = '{98.5699788203};
test_output[1975] = '{3.52940762513e-05};
############ END DEBUG ############*/
test_input[15808:15815] = '{32'hc2af6296, 32'hc14ec887, 32'hc0b3d578, 32'hc11aa4c8, 32'hc0528750, 32'hc27610da, 32'h42022643, 32'h424755c6};
test_label[1976] = '{32'h424755c6};
test_output[1976] = '{32'h330432fe};
/*############ DEBUG ############
test_input[15808:15815] = '{-87.6925488303, -12.9239573018, -5.61980812284, -9.66522973874, -3.28950884736, -61.5164556715, 32.5373642336, 49.8337642063};
test_label[1976] = '{49.8337642063};
test_output[1976] = '{3.07800221163e-08};
############ END DEBUG ############*/
test_input[15816:15823] = '{32'hc28af595, 32'hc207eb1c, 32'hc229d166, 32'h425eacb2, 32'h41e8b5c1, 32'hc29e2f3e, 32'h425ecb21, 32'hc1f3d1ea};
test_label[1977] = '{32'hc1f3d1ea};
test_output[1977] = '{32'h42adb562};
/*############ DEBUG ############
test_input[15816:15823] = '{-69.4796547404, -33.9795995986, -42.4544889146, 55.6686474619, 29.0887472547, -79.0922691392, 55.6983683987, -30.4774966957};
test_label[1977] = '{-30.4774966957};
test_output[1977] = '{86.8542622192};
############ END DEBUG ############*/
test_input[15824:15831] = '{32'hc1e63e84, 32'hc29c0d60, 32'hc2838f2a, 32'h426937ae, 32'hc078c4bf, 32'h422b32cc, 32'h40b27f3b, 32'h410948f1};
test_label[1978] = '{32'hc29c0d60};
test_output[1978] = '{32'h4308549c};
/*############ DEBUG ############
test_input[15824:15831] = '{-28.7805245605, -78.0261217499, -65.7796141394, 58.304376226, -3.88700847706, 42.7996072046, 5.57803092517, 8.58030748634};
test_label[1978] = '{-78.0261217499};
test_output[1978] = '{136.330498161};
############ END DEBUG ############*/
test_input[15832:15839] = '{32'h42695d12, 32'h423a8665, 32'h429d0ded, 32'hc1d0ee3c, 32'h42852f68, 32'hc18f8e8b, 32'hc17d61e5, 32'h3f833084};
test_label[1979] = '{32'h42852f68};
test_output[1979] = '{32'h413ef42e};
/*############ DEBUG ############
test_input[15832:15839] = '{58.3408896758, 46.6312462363, 78.5272008654, -26.1163262893, 66.5925933431, -17.9446019338, -15.8363997797, 1.0249180709};
test_label[1979] = '{66.5925933431};
test_output[1979] = '{11.9346140834};
############ END DEBUG ############*/
test_input[15840:15847] = '{32'h42b84bed, 32'hc24b9ddd, 32'hc2bdb4fa, 32'hc1f599d5, 32'h423610e9, 32'hc230c753, 32'hc2893998, 32'hc29b3bf4};
test_label[1980] = '{32'hc1f599d5};
test_output[1980] = '{32'h42f5b262};
/*############ DEBUG ############
test_input[15840:15847] = '{92.1482901464, -50.9041633346, -94.8534674256, -30.7001133519, 45.5165148861, -44.1946534496, -68.6124900412, -77.6170937206};
test_label[1980] = '{-30.7001133519};
test_output[1980] = '{122.848403498};
############ END DEBUG ############*/
test_input[15848:15855] = '{32'h42baf3ed, 32'hc1a1445f, 32'hc23905b5, 32'hc23e4a06, 32'hc2105dfc, 32'hc220cc53, 32'h420be594, 32'h4285733b};
test_label[1981] = '{32'hc2105dfc};
test_output[1981] = '{32'h43019176};
/*############ DEBUG ############
test_input[15848:15855] = '{93.476419804, -20.1583836673, -46.255573487, -47.5722889833, -36.0917817134, -40.1995359101, 34.9741981145, 66.7250616995};
test_label[1981] = '{-36.0917817134};
test_output[1981] = '{129.568201517};
############ END DEBUG ############*/
test_input[15856:15863] = '{32'hc2b03d55, 32'hc1789316, 32'h41fd0fdc, 32'h429c1243, 32'hc2a3bf46, 32'h420d254c, 32'hc24d0981, 32'h41f891e7};
test_label[1982] = '{32'hc2a3bf46};
test_output[1982] = '{32'h431fe8c5};
/*############ DEBUG ############
test_input[15856:15863] = '{-88.1197889804, -15.5359093977, 31.632743549, 78.0356684688, -81.8735807164, 35.2864209839, -51.2592803076, 31.0712407744};
test_label[1982] = '{-81.8735807164};
test_output[1982] = '{159.909249185};
############ END DEBUG ############*/
test_input[15864:15871] = '{32'h424ac37a, 32'h40831da2, 32'hc2c44211, 32'h42990f4a, 32'hc2c5a9e2, 32'h429850d0, 32'h4000f017, 32'hc210a433};
test_label[1983] = '{32'hc2c5a9e2};
test_output[1983] = '{32'h432fe2d1};
/*############ DEBUG ############
test_input[15864:15871] = '{50.6908935243, 4.09736705414, -98.1290373257, 76.5298593472, -98.8317987164, 76.1578360157, 2.01465392863, -36.1603516937};
test_label[1983] = '{-98.8317987164};
test_output[1983] = '{175.885994894};
############ END DEBUG ############*/
test_input[15872:15879] = '{32'h427ce0f9, 32'hc2b69c23, 32'h424d21e1, 32'hc264d28a, 32'h428f95bf, 32'h409b10b4, 32'h42c3f984, 32'hc29388c0};
test_label[1984] = '{32'h409b10b4};
test_output[1984] = '{32'h42ba4879};
/*############ DEBUG ############
test_input[15872:15879] = '{63.219699017, -91.3049574879, 51.2830835081, -57.2056059253, 71.7924707624, 4.84578872709, 97.9873365783, -73.7670911757};
test_label[1984] = '{4.84578872709};
test_output[1984] = '{93.1415478512};
############ END DEBUG ############*/
test_input[15880:15887] = '{32'h42184d7b, 32'h421ef652, 32'hc2115a4f, 32'h4298f13f, 32'h4281da81, 32'hc223dafb, 32'h426afdad, 32'h42a547ab};
test_label[1985] = '{32'h426afdad};
test_output[1985] = '{32'h41bf2799};
/*############ DEBUG ############
test_input[15880:15887] = '{38.0756646264, 39.7405487391, -36.3381907873, 76.4711809446, 64.9267634945, -40.9638484577, 58.7477319464, 82.6399760769};
test_label[1985] = '{58.7477319464};
test_output[1985] = '{23.8943357191};
############ END DEBUG ############*/
test_input[15888:15895] = '{32'h426d0ec1, 32'h4183b777, 32'h42a079f6, 32'h427d67fb, 32'hc2009e7c, 32'hc1a8543d, 32'h429edaf6, 32'h42a4ae02};
test_label[1986] = '{32'h4183b777};
test_output[1986] = '{32'h42841369};
/*############ DEBUG ############
test_input[15888:15895] = '{59.2644063748, 16.4645827531, 80.2382022144, 63.351542142, -32.1547709404, -21.0411313741, 79.4276608967, 82.3398582562};
test_label[1986] = '{16.4645827531};
test_output[1986] = '{66.0379128978};
############ END DEBUG ############*/
test_input[15896:15903] = '{32'h42b45f15, 32'h42a788d4, 32'h41a3353e, 32'h427485e8, 32'hc198241a, 32'hc13eb187, 32'h41c42cad, 32'hc20cfff9};
test_label[1987] = '{32'h41a3353e};
test_output[1987] = '{32'h428b929b};
/*############ DEBUG ############
test_input[15896:15903] = '{90.1857067005, 83.7672390595, 20.4009965133, 61.130767459, -19.0176268634, -11.9183418202, 24.5218135042, -35.2499730379};
test_label[1987] = '{20.4009965133};
test_output[1987] = '{69.7863400122};
############ END DEBUG ############*/
test_input[15904:15911] = '{32'hc28db630, 32'h429427e7, 32'h40b77b22, 32'hc27a5e12, 32'h42c22f84, 32'hc1faec58, 32'hc2195977, 32'hc16122c3};
test_label[1988] = '{32'h429427e7};
test_output[1988] = '{32'h41b81e74};
/*############ DEBUG ############
test_input[15904:15911] = '{-70.8558329888, 74.0779362039, 5.73378081228, -62.5918643236, 97.0928059459, -31.3654029462, -38.3373683486, -14.0709865901};
test_label[1988] = '{74.0779362039};
test_output[1988] = '{23.0148697421};
############ END DEBUG ############*/
test_input[15912:15919] = '{32'hc1abd73f, 32'hc2a9a1b0, 32'hc2644e1e, 32'h42ba5db3, 32'h429e37b1, 32'hc20f046d, 32'hc293b43f, 32'hc2703cfb};
test_label[1989] = '{32'h42ba5db3};
test_output[1989] = '{32'h354f3df5};
/*############ DEBUG ############
test_input[15912:15919] = '{-21.4801004337, -84.8157940505, -57.0762855579, 93.1830041558, 79.1087707805, -35.7543207472, -73.8520403013, -60.0595528608};
test_label[1989] = '{93.1830041558};
test_output[1989] = '{7.72036690614e-07};
############ END DEBUG ############*/
test_input[15920:15927] = '{32'h40a43bf9, 32'h4293d05a, 32'hc2a2ff06, 32'hc2446567, 32'hc2b4022e, 32'h427766cc, 32'hc19bc198, 32'hc1a69cd6};
test_label[1990] = '{32'h40a43bf9};
test_output[1990] = '{32'h42898c9b};
/*############ DEBUG ############
test_input[15920:15927] = '{5.13232066403, 73.906936948, -81.4980958647, -49.0990271042, -90.0042569753, 61.8503862099, -19.4695278515, -20.8265793999};
test_label[1990] = '{5.13232066403};
test_output[1990] = '{68.7746220903};
############ END DEBUG ############*/
test_input[15928:15935] = '{32'hc225c2e8, 32'hc23244bd, 32'h428ebd01, 32'hc199d31f, 32'h428c07d4, 32'h41a57bcc, 32'hc263d13d, 32'hc24a51e4};
test_label[1991] = '{32'hc24a51e4};
test_output[1991] = '{32'h42f45b90};
/*############ DEBUG ############
test_input[15928:15935] = '{-41.4403384655, -44.5671254442, 71.3691480636, -19.2280858618, 70.0152882181, 20.6854483321, -56.9543327929, -50.5799702378};
test_label[1991] = '{-50.5799702378};
test_output[1991] = '{122.178833462};
############ END DEBUG ############*/
test_input[15936:15943] = '{32'h4162cd63, 32'hc2278005, 32'h423d8eed, 32'hc1b6b488, 32'h4107e376, 32'hc2073389, 32'h427cb92f, 32'h42b22cad};
test_label[1992] = '{32'hc2073389};
test_output[1992] = '{32'h42f5c671};
/*############ DEBUG ############
test_input[15936:15943] = '{14.1751434965, -41.8750180027, 47.3895770739, -22.838150118, 8.49303239577, -33.8003254767, 63.1808452125, 89.0872582769};
test_label[1992] = '{-33.8003254767};
test_output[1992] = '{122.887583754};
############ END DEBUG ############*/
test_input[15944:15951] = '{32'h429d6634, 32'hc16ca7de, 32'hc2a62363, 32'h410c2ac9, 32'hc2a46c82, 32'hc255d604, 32'hc268ce23, 32'h42ace146};
test_label[1993] = '{32'h429d6634};
test_output[1993] = '{32'h40f7b4ab};
/*############ DEBUG ############
test_input[15944:15951] = '{78.6996186054, -14.7909835273, -83.0691175674, 8.76044562293, -82.2119313839, -53.4589986056, -58.2013061154, 86.4399880762};
test_label[1993] = '{78.6996186054};
test_output[1993] = '{7.74080428717};
############ END DEBUG ############*/
test_input[15952:15959] = '{32'h42b6496d, 32'hc1d086dc, 32'hc10483ff, 32'h41f7c595, 32'h41fa1b7a, 32'hc28722c8, 32'h42bd9b53, 32'hc2a37dd6};
test_label[1994] = '{32'h42b6496d};
test_output[1994] = '{32'h406bdd15};
/*############ DEBUG ############
test_input[15952:15959] = '{91.1434076135, -26.065849656, -8.28222552412, 30.9714757342, 31.2634166469, -67.5679290678, 94.803368368, -81.7457746501};
test_label[1994] = '{91.1434076135};
test_output[1994] = '{3.68536874291};
############ END DEBUG ############*/
test_input[15960:15967] = '{32'h42bcb2ae, 32'hc2822306, 32'hc240c36d, 32'hc2225410, 32'hc2a772c2, 32'hc1a89c29, 32'hc268493f, 32'h42a33cfd};
test_label[1995] = '{32'hc268493f};
test_output[1995] = '{32'h43186ba7};
/*############ DEBUG ############
test_input[15960:15967] = '{94.3489832847, -65.068404223, -48.1908445099, -40.5820927001, -83.7241330063, -21.0762492688, -58.0715281417, 81.619116289};
test_label[1995] = '{-58.0715281417};
test_output[1995] = '{152.420514388};
############ END DEBUG ############*/
test_input[15968:15975] = '{32'h423ca54e, 32'h41933d22, 32'h416e6cda, 32'hc1847e2a, 32'hc19c7d7e, 32'h41d083d6, 32'h40f67d42, 32'hc164edc9};
test_label[1996] = '{32'h41933d22};
test_output[1996] = '{32'h41e60d7a};
/*############ DEBUG ############
test_input[15968:15975] = '{47.1614294488, 18.4048491089, 14.9015755225, -16.5616032057, -19.5612762821, 26.0643723994, 7.70279034351, -14.3080525921};
test_label[1996] = '{18.4048491089};
test_output[1996] = '{28.7565803405};
############ END DEBUG ############*/
test_input[15976:15983] = '{32'h424d667d, 32'hc25ff50e, 32'hc294dc35, 32'h42c4acf7, 32'hc24f2c6a, 32'h42b242d4, 32'h42c34d64, 32'h41ccdc30};
test_label[1997] = '{32'hc294dc35};
test_output[1997] = '{32'h432d2cf5};
/*############ DEBUG ############
test_input[15976:15983] = '{51.3500860662, -55.9893129767, -74.4300914906, 98.3378191989, -51.7933719194, 89.1305235358, 97.651156952, 25.6075129607};
test_label[1997] = '{-74.4300914906};
test_output[1997] = '{173.175608841};
############ END DEBUG ############*/
test_input[15984:15991] = '{32'hc199bb7e, 32'hc2242ee9, 32'h41fdf4c3, 32'h4296e100, 32'hc2221c1f, 32'hc235db26, 32'h428d201b, 32'h425769ae};
test_label[1998] = '{32'h41fdf4c3};
test_output[1998] = '{32'h422ecf65};
/*############ DEBUG ############
test_input[15984:15991] = '{-19.2165482034, -41.0458095975, 31.7445121862, 75.4394546365, -40.5274618112, -45.4640119309, 70.5627095192, 53.8532012218};
test_label[1998] = '{31.7445121862};
test_output[1998] = '{43.7025353334};
############ END DEBUG ############*/
test_input[15992:15999] = '{32'hc2686883, 32'hc238722b, 32'hc2bf9400, 32'hc22355f6, 32'hc11ea04c, 32'h42a350ce, 32'h42658fc1, 32'hc191a58d};
test_label[1999] = '{32'hc22355f6};
test_output[1999] = '{32'h42f4fbc9};
/*############ DEBUG ############
test_input[15992:15999] = '{-58.1020636877, -46.1114935945, -95.7890636455, -40.8339472509, -9.91413526301, 81.6578226239, 57.3903848854, -18.2058361081};
test_label[1999] = '{-40.8339472509};
test_output[1999] = '{122.491769875};
############ END DEBUG ############*/
test_input[16000:16007] = '{32'hc1fd7f6e, 32'hbc77a408, 32'hc19bc7ef, 32'hc1f922a6, 32'hc2c32cdb, 32'h42c2d791, 32'hc283c377, 32'h422c89a4};
test_label[2000] = '{32'hc283c377};
test_output[2000] = '{32'h43234d84};
/*############ DEBUG ############
test_input[16000:16007] = '{-31.6872215581, -0.0151147919662, -19.4726246998, -31.141917831, -97.587604783, 97.4210301228, -65.881765173, 43.1344144718};
test_label[2000] = '{-65.881765173};
test_output[2000] = '{163.302795296};
############ END DEBUG ############*/
test_input[16008:16015] = '{32'hc23ea083, 32'h42881c48, 32'h42bb3274, 32'hc256daff, 32'h41833acb, 32'hc247f52d, 32'hc294d967, 32'hc22482e3};
test_label[2001] = '{32'h41833acb};
test_output[2001] = '{32'h429a63c2};
/*############ DEBUG ############
test_input[16008:16015] = '{-47.656748803, 68.0552393019, 93.5985429488, -53.7138616488, 16.4037066478, -49.9894309739, -74.4246163492, -41.1278173205};
test_label[2001] = '{16.4037066478};
test_output[2001] = '{77.194836301};
############ END DEBUG ############*/
test_input[16016:16023] = '{32'hc1847476, 32'h423d237c, 32'h41984dfd, 32'hc23d6324, 32'h417334c9, 32'h427fc1c1, 32'hc2947fb3, 32'hc21d4640};
test_label[2002] = '{32'h417334c9};
test_output[2002] = '{32'h4242f48e};
/*############ DEBUG ############
test_input[16016:16023] = '{-16.5568653921, 47.2846528555, 19.0380794133, -47.3468177814, 15.2003872622, 63.9392116744, -74.2494146336, -39.3186036755};
test_label[2002] = '{15.2003872622};
test_output[2002] = '{48.7388244707};
############ END DEBUG ############*/
test_input[16024:16031] = '{32'h42c73c09, 32'hc265aa25, 32'hc280613e, 32'h41a49a3e, 32'hc23b6e23, 32'hc27c43c8, 32'hc220f576, 32'h421d68cc};
test_label[2003] = '{32'h41a49a3e};
test_output[2003] = '{32'h429e1579};
/*############ DEBUG ############
test_input[16024:16031] = '{99.6172524002, -57.4161566837, -64.1899238957, 20.5753133541, -46.8575569097, -63.0661936313, -40.2397075111, 39.3523401397};
test_label[2003] = '{20.5753133541};
test_output[2003] = '{79.0419390461};
############ END DEBUG ############*/
test_input[16032:16039] = '{32'h42675832, 32'h42c0a46f, 32'hc2388529, 32'h4296a0f1, 32'h42b969ff, 32'hc2a397d1, 32'h42484303, 32'hc22178e5};
test_label[2004] = '{32'h4296a0f1};
test_output[2004] = '{32'h41a8446a};
/*############ DEBUG ############
test_input[16032:16039] = '{57.8361290433, 96.3211613208, -46.1300383923, 75.3143398994, 92.7070245146, -81.7965179018, 50.0654405058, -40.3680591997};
test_label[2004] = '{75.3143398994};
test_output[2004] = '{21.0334050942};
############ END DEBUG ############*/
test_input[16040:16047] = '{32'hbf96626c, 32'h4275fd7d, 32'h42596bec, 32'hc2b31e52, 32'hc1a56392, 32'hc2aff73b, 32'h426d0eb7, 32'h42ae6f3e};
test_label[2005] = '{32'hbf96626c};
test_output[2005] = '{32'h42b0c8c7};
/*############ DEBUG ############
test_input[16040:16047] = '{-1.17487860307, 61.4975477975, 54.3553939232, -89.5592210801, -20.673618022, -87.9828714238, 59.2643689547, 87.2172681658};
test_label[2005] = '{-1.17487860307};
test_output[2005] = '{88.3921467689};
############ END DEBUG ############*/
test_input[16048:16055] = '{32'h42a0ab3a, 32'hc1d0b0b1, 32'h42aea44c, 32'h414a79c3, 32'hc045b6ac, 32'h427462e9, 32'hc22de3ca, 32'hbf1e32e4};
test_label[2006] = '{32'hc22de3ca};
test_output[2006] = '{32'h4302cb55};
/*############ DEBUG ############
test_input[16048:16055] = '{80.3344261723, -26.0862746512, 87.3208919924, 12.6547268331, -3.08927442553, 61.09659081, -43.4724497554, -0.617964026678};
test_label[2006] = '{-43.4724497554};
test_output[2006] = '{130.794265628};
############ END DEBUG ############*/
test_input[16056:16063] = '{32'hc2a18a40, 32'hc2b39e10, 32'h423bf5b8, 32'hc251b36b, 32'h4299f715, 32'h41cb97fd, 32'h422a4774, 32'hc2866ea8};
test_label[2007] = '{32'hc2a18a40};
test_output[2007] = '{32'h431dc0aa};
/*############ DEBUG ############
test_input[16056:16063] = '{-80.7700175553, -89.8087158905, 46.9899604079, -52.4252128935, 76.9825838392, 25.4492134171, 42.5697802316, -67.2161239429};
test_label[2007] = '{-80.7700175553};
test_output[2007] = '{157.752601395};
############ END DEBUG ############*/
test_input[16064:16071] = '{32'h404a7508, 32'hc2bdfc11, 32'h4182a102, 32'h4249cd27, 32'hc13ac6da, 32'h42057182, 32'hc22c4855, 32'h40164040};
test_label[2008] = '{32'hc22c4855};
test_output[2008] = '{32'h42bb0abe};
/*############ DEBUG ############
test_input[16064:16071] = '{3.16339293308, -94.9923159607, 16.3286174118, 50.4503434733, -11.6735474201, 33.3608481733, -43.0706350808, 2.34767162525};
test_label[2008] = '{-43.0706350808};
test_output[2008] = '{93.5209785919};
############ END DEBUG ############*/
test_input[16072:16079] = '{32'h4199dfa8, 32'h428cd0f6, 32'h42bf8e25, 32'h4211920a, 32'hc20e0408, 32'h422cb923, 32'h40aa81a5, 32'hc1d44f67};
test_label[2009] = '{32'hc20e0408};
test_output[2009] = '{32'h43034814};
/*############ DEBUG ############
test_input[16072:16079] = '{19.2342076425, 70.4081238074, 95.7776238457, 36.3926159891, -35.5039377164, 43.1807968412, 5.32832592687, -26.5387712357};
test_label[2009] = '{-35.5039377164};
test_output[2009] = '{131.281561562};
############ END DEBUG ############*/
test_input[16080:16087] = '{32'hc2aab5de, 32'hc28c4196, 32'h424fce6d, 32'hc29e8fed, 32'hc0ef14f3, 32'hc263c4ce, 32'hc2a88fa1, 32'h3e2bbe37};
test_label[2010] = '{32'hc0ef14f3};
test_output[2010] = '{32'h426db10c};
/*############ DEBUG ############
test_input[16080:16087] = '{-85.3552070417, -70.1280973607, 51.9515890371, -79.2811028632, -7.47130736868, -56.9421922296, -84.2805264242, 0.167717798721};
test_label[2010] = '{-7.47130736868};
test_output[2010] = '{59.4228964058};
############ END DEBUG ############*/
test_input[16088:16095] = '{32'hc21a2641, 32'h42185f1f, 32'hc1d86c78, 32'h41a379ba, 32'hc17f9199, 32'hc206c54b, 32'hc2947940, 32'h422f1e4f};
test_label[2011] = '{32'hc206c54b};
test_output[2011] = '{32'h429af389};
/*############ DEBUG ############
test_input[16088:16095] = '{-38.5373558336, 38.0928908605, -27.0529641951, 20.4344370209, -15.9730460173, -33.6926672988, -74.2368136329, 43.7795997812};
test_label[2011] = '{-33.6926672988};
test_output[2011] = '{77.4756520783};
############ END DEBUG ############*/
test_input[16096:16103] = '{32'h423b092a, 32'h42a08bf5, 32'hc29bba0e, 32'h422e588e, 32'h422c55f6, 32'h40eeb351, 32'h41cc574a, 32'hc2af89ff};
test_label[2012] = '{32'h423b092a};
test_output[2012] = '{32'h42060ec0};
/*############ DEBUG ############
test_input[16096:16103] = '{46.758949536, 80.2733539351, -77.8633850772, 43.5864774434, 43.0839443537, 7.45938942786, 25.5426209471, -87.7695268903};
test_label[2012] = '{46.758949536};
test_output[2012] = '{33.5144043991};
############ END DEBUG ############*/
test_input[16104:16111] = '{32'hc1d16ad9, 32'hc2938b5c, 32'h42815777, 32'hc2a36163, 32'h41a7f1cc, 32'h42b643cb, 32'h4230dc48, 32'hc2ba705d};
test_label[2013] = '{32'h41a7f1cc};
test_output[2013] = '{32'h428c4758};
/*############ DEBUG ############
test_input[16104:16111] = '{-26.1771717409, -73.7721866233, 64.6708287907, -81.6902110973, 20.9930644463, 91.1324105312, 44.215118032, -93.219461331};
test_label[2013] = '{20.9930644463};
test_output[2013] = '{70.1393460849};
############ END DEBUG ############*/
test_input[16112:16119] = '{32'h42771a9a, 32'h4220a526, 32'hc13972c3, 32'hc21801a5, 32'h42a78780, 32'h42c0f5d3, 32'h40142ed5, 32'h421dc447};
test_label[2014] = '{32'h42c0f5d3};
test_output[2014] = '{32'h36499ca7};
/*############ DEBUG ############
test_input[16112:16119] = '{61.7759788991, 40.1612777046, -11.5905178035, -38.0016057477, 83.7646457349, 96.4801262461, 2.31535846496, 39.4416788869};
test_label[2014] = '{96.4801262461};
test_output[2014] = '{3.00425177872e-06};
############ END DEBUG ############*/
test_input[16120:16127] = '{32'hc0696df1, 32'hc1adc042, 32'h41990125, 32'hc2060cfc, 32'hc2323215, 32'h4285ea2c, 32'hc24c6287, 32'h41ff314e};
test_label[2015] = '{32'h4285ea2c};
test_output[2015] = '{32'h26200000};
/*############ DEBUG ############
test_input[16120:16127] = '{-3.64733533104, -21.7188752465, 19.1255596154, -33.512681774, -44.5489100896, 66.9573661671, -51.0962173345, 31.8990742987};
test_label[2015] = '{66.9573661671};
test_output[2015] = '{5.55111512313e-16};
############ END DEBUG ############*/
test_input[16128:16135] = '{32'hc2629c91, 32'h42a6b95c, 32'hc18c5833, 32'h4279e66d, 32'hc0b9d1d0, 32'h40ecaadd, 32'h429d047d, 32'hc2a38d82};
test_label[2016] = '{32'hc0b9d1d0};
test_output[2016] = '{32'h42b25a74};
/*############ DEBUG ############
test_input[16128:16135] = '{-56.6528979601, 83.3620315444, -17.5430664378, 62.4750251665, -5.80686174131, 7.39585743251, 78.5087647794, -81.7763854066};
test_label[2016] = '{-5.80686174131};
test_output[2016] = '{89.1766658475};
############ END DEBUG ############*/
test_input[16136:16143] = '{32'h4246ecf4, 32'hc2074256, 32'hc1035941, 32'h423327d8, 32'h4232780f, 32'hc2960baa, 32'h417407e3, 32'hc2b0a672};
test_label[2017] = '{32'hc1035941};
test_output[2017] = '{32'h4267d0a4};
/*############ DEBUG ############
test_input[16136:16143] = '{49.7313987376, -33.8147802579, -8.20929056014, 44.7889083669, 44.6172454051, -75.0227830211, 15.2519258453, -88.3250856806};
test_label[2017] = '{-8.20929056014};
test_output[2017] = '{57.9537514828};
############ END DEBUG ############*/
test_input[16144:16151] = '{32'h42094b49, 32'hc118eb7b, 32'h423f5b32, 32'h410d9f86, 32'hc2af8915, 32'hc244e854, 32'h422dd3a6, 32'h425cec34};
test_label[2018] = '{32'h42094b49};
test_output[2018] = '{32'h41a7431d};
/*############ DEBUG ############
test_input[16144:16151] = '{34.3235219881, -9.557490415, 47.839056587, 8.85144638971, -87.7677412586, -49.2268834835, 43.45668899, 55.2306678008};
test_label[2018] = '{34.3235219881};
test_output[2018] = '{20.9077697232};
############ END DEBUG ############*/
test_input[16152:16159] = '{32'hc12f7842, 32'hc2767981, 32'h4163f531, 32'hc2170458, 32'h41b514bc, 32'hc2500ef7, 32'hc2894e27, 32'h42b114ff};
test_label[2019] = '{32'hc2767981};
test_output[2019] = '{32'h431628e0};
/*############ DEBUG ############
test_input[16152:16159] = '{-10.9668595663, -61.6186544662, 14.2473611193, -37.7542410967, 22.6351245806, -52.014613836, -68.6526429188, 88.5410099441};
test_label[2019] = '{-61.6186544662};
test_output[2019] = '{150.15966441};
############ END DEBUG ############*/
test_input[16160:16167] = '{32'hc259bfeb, 32'h4294a001, 32'hc283a4ee, 32'h4291f26b, 32'h4123a2b3, 32'hc2b1d0ac, 32'h423adb07, 32'hc2bb6246};
test_label[2020] = '{32'hc283a4ee};
test_output[2020] = '{32'h430c5e0f};
/*############ DEBUG ############
test_input[16160:16167] = '{-54.437420828, 74.312509588, -65.8221301223, 72.9734690147, 10.227221532, -88.9075591182, 46.713892148, -93.6919437728};
test_label[2020] = '{-65.8221301223};
test_output[2020] = '{140.367414342};
############ END DEBUG ############*/
test_input[16168:16175] = '{32'hc1fbfaea, 32'h425b3967, 32'h429a73c3, 32'h41f12cdb, 32'h42bc2fae, 32'hc24a3077, 32'hc160a2fb, 32'h42a5a5fa};
test_label[2021] = '{32'h429a73c3};
test_output[2021] = '{32'h4186efb4};
/*############ DEBUG ############
test_input[16168:16175] = '{-31.4975157602, 54.8060554071, 77.226095812, 30.1469026836, 94.0931257253, -50.5473296783, -14.0397896808, 82.8241735827};
test_label[2021] = '{77.226095812};
test_output[2021] = '{16.8670427237};
############ END DEBUG ############*/
test_input[16176:16183] = '{32'hc1638271, 32'h420f75f4, 32'h40f45e0f, 32'h42a3c90f, 32'hc2aa442e, 32'h42c5a2e3, 32'hc1bb6cc8, 32'hc1f2a944};
test_label[2022] = '{32'hc1638271};
test_output[2022] = '{32'h42e21331};
/*############ DEBUG ############
test_input[16176:16183] = '{-14.2193460885, 35.8651896848, 7.63648170556, 81.8926915481, -85.1331598531, 98.8181378065, -23.4281160893, -30.332649698};
test_label[2022] = '{-14.2193460885};
test_output[2022] = '{113.03748394};
############ END DEBUG ############*/
test_input[16184:16191] = '{32'h423efb49, 32'h42420efb, 32'hc2671d3e, 32'h427803d9, 32'hc25555d0, 32'h425a8873, 32'h415996c5, 32'h4195ffb4};
test_label[2023] = '{32'h4195ffb4};
test_output[2023] = '{32'h422d04a4};
/*############ DEBUG ############
test_input[16184:16191] = '{47.7453939557, 48.5146312441, -57.7785572271, 62.0037563549, -53.3338023243, 54.6332509657, 13.5993087692, 18.7498558275};
test_label[2023] = '{18.7498558275};
test_output[2023] = '{43.2545319062};
############ END DEBUG ############*/
test_input[16192:16199] = '{32'hc1845b10, 32'h423e8cea, 32'hc292ba91, 32'h4283aa97, 32'hc1271cd7, 32'hc2338172, 32'h4282d4b4, 32'h41b64c81};
test_label[2024] = '{32'hc1845b10};
test_output[2024] = '{32'h42a5c464};
/*############ DEBUG ############
test_input[16192:16199] = '{-16.5444632391, 47.6376102357, -73.3643887104, 65.833185948, -10.4445410603, -44.8764126945, 65.4154353859, 22.7873560461};
test_label[2024] = '{-16.5444632391};
test_output[2024] = '{82.8835787337};
############ END DEBUG ############*/
test_input[16200:16207] = '{32'hc1dde44f, 32'hc2588a34, 32'hc100c01a, 32'hc218a741, 32'h428ad7a5, 32'hc1f8e399, 32'h422ba0fb, 32'hc2341bde};
test_label[2025] = '{32'hc218a741};
test_output[2025] = '{32'h42d72b45};
/*############ DEBUG ############
test_input[16200:16207] = '{-27.7364780617, -54.1349650659, -8.04689982893, -38.1633341423, 69.4211785897, -31.1111322334, 42.9072065972, -45.0272138083};
test_label[2025] = '{-38.1633341423};
test_output[2025] = '{107.584512732};
############ END DEBUG ############*/
test_input[16208:16215] = '{32'h4276262d, 32'h424d19f2, 32'hc2881fd5, 32'h41da87fa, 32'hc297935a, 32'h42681c9e, 32'h412cb97a, 32'hc29edae7};
test_label[2026] = '{32'h41da87fa};
test_output[2026] = '{32'h42090068};
/*############ DEBUG ############
test_input[16208:16215] = '{61.5372818798, 51.2753355771, -68.0621720488, 27.3163953696, -75.7877991076, 58.027948181, 10.7952826336, -79.4275434074};
test_label[2026] = '{27.3163953696};
test_output[2026] = '{34.250398495};
############ END DEBUG ############*/
test_input[16216:16223] = '{32'h412e841c, 32'hc10d1a42, 32'h42a7f49c, 32'h3feb9c86, 32'hc2c644a2, 32'hc1baea80, 32'hc0dec60a, 32'hc2bd4d09};
test_label[2027] = '{32'hc2bd4d09};
test_output[2027] = '{32'h4332a0d3};
/*############ DEBUG ############
test_input[16216:16223] = '{10.9072532911, -8.81891061251, 83.9777564526, 1.84071416406, -99.1340468841, -23.3645013263, -6.96167455875, -94.6504562295};
test_label[2027] = '{-94.6504562295};
test_output[2027] = '{178.628212682};
############ END DEBUG ############*/
test_input[16224:16231] = '{32'h42ac20e4, 32'hc1fc6ebf, 32'hc2273e7f, 32'hc295beb0, 32'h428fa360, 32'hc184f324, 32'h426ed00f, 32'h42879b4f};
test_label[2028] = '{32'hc295beb0};
test_output[2028] = '{32'h4320efca};
/*############ DEBUG ############
test_input[16224:16231] = '{86.0642373442, -31.554076075, -41.8110320044, -74.872435915, 71.8190955877, -16.6187213778, 59.7031840389, 67.8033389714};
test_label[2028] = '{-74.872435915};
test_output[2028] = '{160.936673922};
############ END DEBUG ############*/
test_input[16232:16239] = '{32'hc2c3fa2b, 32'hc0fee484, 32'h428bc0c2, 32'h42082bc1, 32'h418deb73, 32'h42b6f071, 32'hc0e0ba19, 32'hc11e7bef};
test_label[2029] = '{32'hc2c3fa2b};
test_output[2029] = '{32'h433d754e};
/*############ DEBUG ############
test_input[16232:16239] = '{-97.9886097686, -7.96539492567, 69.8764777355, 34.0427276232, 17.7399657489, 91.4696090315, -7.02271711738, -9.90525760797};
test_label[2029] = '{-97.9886097686};
test_output[2029] = '{189.4582188};
############ END DEBUG ############*/
test_input[16240:16247] = '{32'hc1a10c48, 32'hc2365500, 32'hc23d3265, 32'h42900963, 32'h41906fec, 32'h3b655190, 32'hc2012e52, 32'h4261a06c};
test_label[2030] = '{32'h3b655190};
test_output[2030] = '{32'h42900799};
/*############ DEBUG ############
test_input[16240:16247] = '{-20.1309971879, -45.5830066864, -47.299212131, 72.0183355905, 18.0546491137, 0.0034991241032, -32.2952336697, 56.4066632101};
test_label[2030] = '{0.0034991241032};
test_output[2030] = '{72.0148366323};
############ END DEBUG ############*/
test_input[16248:16255] = '{32'hc273e022, 32'h4233bc84, 32'hc2becae9, 32'hc2ab2507, 32'h42bf3f28, 32'hc23a7070, 32'h412f4eeb, 32'h40741930};
test_label[2031] = '{32'h40741930};
test_output[2031] = '{32'h42b79e5e};
/*############ DEBUG ############
test_input[16248:16255] = '{-60.9688786516, 44.9340991743, -95.3963113172, -85.5723193805, 95.6233490998, -46.6098037869, 10.9567666781, 3.81403743262};
test_label[2031] = '{3.81403743262};
test_output[2031] = '{91.8093116672};
############ END DEBUG ############*/
test_input[16256:16263] = '{32'h429fb937, 32'hc21329c7, 32'h4213ca69, 32'hc1b7854e, 32'h412c8590, 32'h41d8b43f, 32'hc22e28f1, 32'hc28ff9ca};
test_label[2032] = '{32'h4213ca69};
test_output[2032] = '{32'h422ba804};
/*############ DEBUG ############
test_input[16256:16263] = '{79.8617455855, -36.7907965729, 36.9476674043, -22.9400897412, 10.782607956, 27.0880113252, -43.5399826917, -71.9878690644};
test_label[2032] = '{36.9476674043};
test_output[2032] = '{42.9140781812};
############ END DEBUG ############*/
test_input[16264:16271] = '{32'h42513c08, 32'h3fc4a1a0, 32'hc292d49f, 32'hc2baf97a, 32'h4266a59d, 32'hc20959d1, 32'h41a59086, 32'hc2a2d2c9};
test_label[2033] = '{32'h41a59086};
test_output[2033] = '{32'h4213e22f};
/*############ DEBUG ############
test_input[16264:16271] = '{52.3086244879, 1.53618239958, -73.4152766305, -93.4872600871, 57.6617302279, -34.3377107358, 20.6955686251, -81.4116895305};
test_label[2033] = '{20.6955686251};
test_output[2033] = '{36.9708838627};
############ END DEBUG ############*/
test_input[16272:16279] = '{32'hc27354d1, 32'h429f0a2c, 32'hc2a7dca2, 32'hc28e6163, 32'h4227bfdc, 32'hc1d6bc48, 32'hc28b5931, 32'hc243f7c9};
test_label[2034] = '{32'h4227bfdc};
test_output[2034] = '{32'h4216547b};
/*############ DEBUG ############
test_input[16272:16279] = '{-60.8328275454, 79.5198634549, -83.9309212318, -71.190206129, 41.9373616863, -26.8419338586, -69.6742042992, -48.991978979};
test_label[2034] = '{41.9373616863};
test_output[2034] = '{37.5825017685};
############ END DEBUG ############*/
test_input[16280:16287] = '{32'hc0937d9f, 32'h4251a21d, 32'hc02e337f, 32'hc2b04227, 32'hc22240e6, 32'hc13ba966, 32'h42102f9a, 32'h42541e4f};
test_label[2035] = '{32'h4251a21d};
test_output[2035] = '{32'h3f869065};
/*############ DEBUG ############
test_input[16280:16287] = '{-4.60908471113, 52.4083131457, -2.72189309241, -88.1292057481, -40.5633758374, -11.7288572395, 36.0464842273, 53.029596791};
test_label[2035] = '{52.4083131457};
test_output[2035] = '{1.05128160875};
############ END DEBUG ############*/
test_input[16288:16295] = '{32'hc2b931e6, 32'hc1157120, 32'hc2c02e71, 32'hc105a216, 32'hc1d1790f, 32'hc2572757, 32'h424f8269, 32'h42827276};
test_label[2036] = '{32'hc2c02e71};
test_output[2036] = '{32'h43215074};
/*############ DEBUG ############
test_input[16288:16295] = '{-92.5974547805, -9.34011797954, -96.0907081314, -8.35207186689, -26.1841106914, -53.7884161734, 51.8773538467, 65.2235576637};
test_label[2036] = '{-96.0907081314};
test_output[2036] = '{161.314267394};
############ END DEBUG ############*/
test_input[16296:16303] = '{32'hc269087e, 32'h42a42e66, 32'hc236e769, 32'h420bb0af, 32'hc1ef316b, 32'h406bd1f0, 32'h4180ba33, 32'h4250737b};
test_label[2037] = '{32'hc236e769};
test_output[2037] = '{32'h42ffa21b};
/*############ DEBUG ############
test_input[16296:16303] = '{-58.2582913572, 82.0906245649, -45.7259848056, 34.9225436736, -29.8991301275, 3.68468859717, 16.0909184342, 52.1127752355};
test_label[2037] = '{-45.7259848056};
test_output[2037] = '{127.81660937};
############ END DEBUG ############*/
test_input[16304:16311] = '{32'hc20fb07f, 32'hc2446522, 32'h4201b35a, 32'hc1aab447, 32'hc2b5e970, 32'hc2903027, 32'h41064a66, 32'h41aa87e4};
test_label[2038] = '{32'hc1aab447};
test_output[2038] = '{32'h42570d81};
/*############ DEBUG ############
test_input[16304:16311] = '{-35.9223579147, -49.09876338, 32.4251483981, -21.3380257612, -90.9559306634, -72.0940479737, 8.39316357932, 21.3163530773};
test_label[2038] = '{-21.3380257612};
test_output[2038] = '{53.7631891392};
############ END DEBUG ############*/
test_input[16312:16319] = '{32'h42471628, 32'hc210c03e, 32'hc2a75860, 32'h429322d4, 32'h423766f4, 32'h4239e1be, 32'hc2b73a53, 32'h416cd5b0};
test_label[2039] = '{32'hc2b73a53};
test_output[2039] = '{32'h43252e93};
/*############ DEBUG ############
test_input[16312:16319] = '{49.7716364652, -36.1877348605, -83.6726076426, 73.5680208067, 45.8505408675, 46.4704508647, -91.613914946, 14.802169353};
test_label[2039] = '{-91.613914946};
test_output[2039] = '{165.181935753};
############ END DEBUG ############*/
test_input[16320:16327] = '{32'h41d3ec81, 32'hc29ba2d2, 32'hc22a4524, 32'h429bc102, 32'hc2b1c1ff, 32'hc23a1c27, 32'hc2884f03, 32'h42031b3e};
test_label[2040] = '{32'hc29ba2d2};
test_output[2040] = '{32'h431bb1ea};
/*############ DEBUG ############
test_input[16320:16327] = '{26.4904803548, -77.8180082226, -42.5675183439, 77.8769669735, -88.8789016747, -46.5274936262, -68.1543226723, 32.7766044379};
test_label[2040] = '{-77.8180082226};
test_output[2040] = '{155.694975196};
############ END DEBUG ############*/
test_input[16328:16335] = '{32'hc16ae6d2, 32'h41b132ca, 32'h42a9664d, 32'hc16949be, 32'h42b2f9af, 32'hc2024a67, 32'hc2138536, 32'h4186a221};
test_label[2041] = '{32'h4186a221};
test_output[2041] = '{32'h42915566};
/*############ DEBUG ############
test_input[16328:16335] = '{-14.6813523956, 22.1497984204, 84.6998056069, -14.580503505, 89.487665368, -32.5726568629, -36.8800890808, 16.8291650503};
test_label[2041] = '{16.8291650503};
test_output[2041] = '{72.6667960796};
############ END DEBUG ############*/
test_input[16336:16343] = '{32'hc2abbc71, 32'hc293bc21, 32'h42626116, 32'hc29e05d2, 32'hc2b53b6e, 32'hc0db4215, 32'h42366046, 32'h42ab97c3};
test_label[2042] = '{32'hc293bc21};
test_output[2042] = '{32'h431fa9f2};
/*############ DEBUG ############
test_input[16336:16343] = '{-85.8680529189, -73.8674366092, 56.594812005, -79.0113676586, -90.6160712259, -6.85181678565, 45.5940175542, 85.7964074864};
test_label[2042] = '{-73.8674366092};
test_output[2042] = '{159.663844096};
############ END DEBUG ############*/
test_input[16344:16351] = '{32'h41a1476d, 32'hc1c98ad0, 32'hc2bd61a9, 32'h42999e8a, 32'hc2a2a99c, 32'h42a51ca2, 32'hc28721bd, 32'hc1b6cd6a};
test_label[2043] = '{32'hc1b6cd6a};
test_output[2043] = '{32'h42d2d19e};
/*############ DEBUG ############
test_input[16344:16351] = '{20.1598754276, -25.1927802926, -94.6907424284, 76.8096479729, -81.3312646387, 82.5559199929, -67.5658955555, -22.850300594};
test_label[2043] = '{-22.850300594};
test_output[2043] = '{105.409410163};
############ END DEBUG ############*/
test_input[16352:16359] = '{32'hc2270cc5, 32'h422048d5, 32'hc2a28eea, 32'h42ad2548, 32'h42abb9a9, 32'hc292a91d, 32'hc1bcb0ed, 32'hc28d28df};
test_label[2044] = '{32'hc2a28eea};
test_output[2044] = '{32'h43284073};
/*############ DEBUG ############
test_input[16352:16359] = '{-41.7624684304, 40.0711232714, -81.2791320731, 86.5728167023, 85.862615541, -73.3303024253, -23.586389494, -70.5798257852};
test_label[2044] = '{-81.2791320731};
test_output[2044] = '{168.251761477};
############ END DEBUG ############*/
test_input[16360:16367] = '{32'h40ed25b6, 32'h42bd15ac, 32'hc282e67b, 32'hc2c488cb, 32'hc271c8ab, 32'hc249e17b, 32'hc23e25b6, 32'hc2c6cac6};
test_label[2045] = '{32'hc249e17b};
test_output[2045] = '{32'h43110334};
/*############ DEBUG ############
test_input[16360:16367] = '{7.41085330842, 94.5423253933, -65.4501591344, -98.2671743801, -60.4459641412, -50.4701943973, -47.5368269509, -99.3960452832};
test_label[2045] = '{-50.4701943973};
test_output[2045] = '{145.012519791};
############ END DEBUG ############*/
test_input[16368:16375] = '{32'hc222debd, 32'hc0c50ce0, 32'h403c2ae3, 32'hc2470f0c, 32'hc1e5719d, 32'hc1efe018, 32'h42a422b5, 32'h41c04212};
test_label[2046] = '{32'hc2470f0c};
test_output[2046] = '{32'h4303d51e};
/*############ DEBUG ############
test_input[16368:16375] = '{-40.7175161498, -6.15782166035, 2.94011763007, -49.7646937019, -28.6804742884, -29.9844199392, 82.0677893591, 24.0322607929};
test_label[2046] = '{-49.7646937019};
test_output[2046] = '{131.832483061};
############ END DEBUG ############*/
test_input[16376:16383] = '{32'h4182aec1, 32'hc28af516, 32'hc2bed121, 32'h429a0297, 32'h42062419, 32'h41dd854e, 32'hc271182c, 32'hc289d3d6};
test_label[2047] = '{32'hc28af516};
test_output[2047] = '{32'h43127bd7};
/*############ DEBUG ############
test_input[16376:16383] = '{16.3353292535, -69.4786837864, -95.4084548957, 77.0050613007, 33.5352526364, 27.6900893893, -60.2736057465, -68.9137431095};
test_label[2047] = '{-69.4786837864};
test_output[2047] = '{146.483745087};
############ END DEBUG ############*/
test_input[16384:16391] = '{32'h42770d89, 32'h41263297, 32'hc1fa65f1, 32'hc212c633, 32'hc2533bf3, 32'hc2b69540, 32'hc26f49ec, 32'h42a85708};
test_label[2048] = '{32'hc2b69540};
test_output[2048] = '{32'h432f7624};
/*############ DEBUG ############
test_input[16384:16391] = '{61.7632194974, 10.387351386, -31.2997759838, -36.693553069, -52.8085423146, -91.2915007638, -59.8221900117, 84.1699819453};
test_label[2048] = '{-91.2915007638};
test_output[2048] = '{175.461482709};
############ END DEBUG ############*/
test_input[16392:16399] = '{32'hc18be064, 32'hc215525c, 32'h42279367, 32'hc2b9d055, 32'hc2628c2c, 32'h42406676, 32'hc1a3e16e, 32'h42bb92cc};
test_label[2049] = '{32'hc2b9d055};
test_output[2049] = '{32'h433ab191};
/*############ DEBUG ############
test_input[16392:16399] = '{-17.484564893, -37.3304295861, 41.8939494505, -92.9068957891, -56.6368861994, 48.1000594137, -20.4850737802, 93.7867156852};
test_label[2049] = '{-92.9068957891};
test_output[2049] = '{186.693611474};
############ END DEBUG ############*/
test_input[16400:16407] = '{32'h42b9e612, 32'hc20b0038, 32'hc119ac59, 32'hc2a188ec, 32'hc1b38752, 32'hc2b5af69, 32'hc2b49535, 32'hc2287ae1};
test_label[2050] = '{32'hc2b49535};
test_output[2050] = '{32'h43373da3};
/*############ DEBUG ############
test_input[16400:16407] = '{92.949352874, -34.7502151842, -9.60457736476, -80.7674284803, -22.4410735909, -90.8425958479, -90.291417094, -42.1199996366};
test_label[2050] = '{-90.291417094};
test_output[2050] = '{183.240769968};
############ END DEBUG ############*/
test_input[16408:16415] = '{32'h42970efb, 32'h417e1f06, 32'h424e88eb, 32'hc1ee3216, 32'hc1f08e09, 32'hc2964a98, 32'h42a6c8db, 32'hc2b7797e};
test_label[2051] = '{32'hc1ee3216};
test_output[2051] = '{32'h42e25593};
/*############ DEBUG ############
test_input[16408:16415] = '{75.5292554872, 15.8825736599, 51.6337074999, -29.774455112, -30.0693525395, -75.145690606, 83.3922940946, -91.737290678};
test_label[2051] = '{-29.774455112};
test_output[2051] = '{113.167133836};
############ END DEBUG ############*/
test_input[16416:16423] = '{32'hc2ab646e, 32'h428ceca7, 32'hc21ee5f5, 32'hc20189be, 32'hc297b1f9, 32'hc20f0d5e, 32'hc25c396c, 32'hc09baa84};
test_label[2052] = '{32'hc2ab646e};
test_output[2052] = '{32'h431c288b};
/*############ DEBUG ############
test_input[16416:16423] = '{-85.6961532466, 70.4622132776, -39.7245660773, -32.3845127432, -75.8476000341, -35.7630548413, -55.0560766134, -4.86456475469};
test_label[2052] = '{-85.6961532466};
test_output[2052] = '{156.158366524};
############ END DEBUG ############*/
test_input[16424:16431] = '{32'hc298f79c, 32'h423436fa, 32'h427b1270, 32'h42122729, 32'hc0e1ed71, 32'h4291c293, 32'hc2515ebc, 32'h410e9825};
test_label[2053] = '{32'hc2515ebc};
test_output[2053] = '{32'h42fa71f7};
/*############ DEBUG ############
test_input[16424:16431] = '{-76.4836103569, 45.0536888725, 62.7680040039, 36.5382414397, -7.06023434691, 72.8800297679, -52.3425147062, 8.91214421387};
test_label[2053] = '{-52.3425147062};
test_output[2053] = '{125.222585062};
############ END DEBUG ############*/
test_input[16432:16439] = '{32'hc04b7072, 32'hc29c9317, 32'hc2927d81, 32'h420882d6, 32'hc2831680, 32'hc2058faf, 32'hc282d641, 32'hc10d1904};
test_label[2054] = '{32'hc04b7072};
test_output[2054] = '{32'h421539dd};
/*############ DEBUG ############
test_input[16432:16439] = '{-3.17873812903, -78.2872858524, -73.2451249667, 34.1277690612, -65.5439471551, -33.3903162819, -65.4184613852, -8.81860718437};
test_label[2054] = '{-3.17873812903};
test_output[2054] = '{37.3065071903};
############ END DEBUG ############*/
test_input[16440:16447] = '{32'h425c3823, 32'hc2c5da52, 32'h4195aa78, 32'h4218a8be, 32'h41cf57a1, 32'h42ac4f13, 32'hc2c359a3, 32'hc13ce014};
test_label[2055] = '{32'h41cf57a1};
test_output[2055] = '{32'h4270f255};
/*############ DEBUG ############
test_input[16440:16447] = '{55.0548202694, -98.9264044676, 18.7082359157, 38.1647857771, 25.9177875114, 86.1544407162, -97.6750726604, -11.8047066067};
test_label[2055] = '{25.9177875114};
test_output[2055] = '{60.2366532048};
############ END DEBUG ############*/
test_input[16448:16455] = '{32'hc182f961, 32'h40ce472c, 32'hc1ebd25c, 32'h412f348a, 32'h4279dfba, 32'hc287ea69, 32'hc1baa0b0, 32'hc168f857};
test_label[2056] = '{32'hc1ebd25c};
test_output[2056] = '{32'h42b7e474};
/*############ DEBUG ############
test_input[16448:16455] = '{-16.3717668304, 6.44618792845, -29.4777154459, 10.9503268514, 62.4684824364, -67.9578299837, -23.3284599761, -14.5606299598};
test_label[2056] = '{-29.4777154459};
test_output[2056] = '{91.9461978823};
############ END DEBUG ############*/
test_input[16456:16463] = '{32'h41be794e, 32'h412a60ba, 32'hc2871945, 32'h42b610df, 32'hc1284087, 32'hc29bba09, 32'h40b29275, 32'h3f9375db};
test_label[2057] = '{32'h3f9375db};
test_output[2057] = '{32'h42b3c308};
/*############ DEBUG ############
test_input[16456:16463] = '{23.8092308231, 10.6486144288, -67.5493522291, 91.0329541991, -10.5157540819, -77.8633488321, 5.58037829201, 1.15203418948};
test_label[2057] = '{1.15203418948};
test_output[2057] = '{89.8809200096};
############ END DEBUG ############*/
test_input[16464:16471] = '{32'hc2a95d59, 32'hc28b6efb, 32'hc298a76a, 32'h422a94ab, 32'h42aeaefa, 32'hc2153970, 32'hc2aff923, 32'h42a4477d};
test_label[2058] = '{32'hc2aff923};
test_output[2058] = '{32'h432f5576};
/*############ DEBUG ############
test_input[16464:16471] = '{-84.6823213697, -69.7167571438, -76.3269842558, 42.6451839633, 87.341747914, -37.306092458, -87.9865938384, 82.1396250936};
test_label[2058] = '{-87.9865938384};
test_output[2058] = '{175.333831522};
############ END DEBUG ############*/
test_input[16472:16479] = '{32'h42090cdf, 32'h42c7911e, 32'h425cc86e, 32'hc21e5eee, 32'hc2c1f32b, 32'hc1d81b9a, 32'hc11f89d2, 32'hc1c46aab};
test_label[2059] = '{32'hc11f89d2};
test_output[2059] = '{32'h42db8258};
/*############ DEBUG ############
test_input[16472:16479] = '{34.2625712389, 99.7834325715, 55.1957327927, -39.5927035178, -96.9749410394, -27.0134772872, -9.97114753934, -24.5520841154};
test_label[2059] = '{-9.97114753934};
test_output[2059] = '{109.754580111};
############ END DEBUG ############*/
test_input[16480:16487] = '{32'h42c0b791, 32'h42ac5f3a, 32'h42c3121f, 32'h4280e7a2, 32'h41774625, 32'h41201f8f, 32'h42806a3e, 32'hc1eebb34};
test_label[2060] = '{32'h42c3121f};
test_output[2060] = '{32'h3e899222};
/*############ DEBUG ############
test_input[16480:16487] = '{96.3585249986, 86.1859916732, 97.5353959981, 64.4524113038, 15.4546255979, 10.0077051407, 64.207501845, -29.8414071382};
test_label[2060] = '{97.5353959981};
test_output[2060] = '{0.268693038711};
############ END DEBUG ############*/
test_input[16488:16495] = '{32'h422a8362, 32'hc2bfaeb4, 32'hc295fdcf, 32'h41791bf2, 32'h3f4e2208, 32'hc16e3b4c, 32'h42909322, 32'h42880cb6};
test_label[2061] = '{32'hc295fdcf};
test_output[2061] = '{32'h43134c0d};
/*############ DEBUG ############
test_input[16488:16495] = '{42.6283046682, -95.8412157087, -74.9957231796, 15.5693229195, 0.805206797814, -14.889476637, 72.2873652927, 68.0248254056};
test_label[2061] = '{-74.9957231796};
test_output[2061] = '{147.297076659};
############ END DEBUG ############*/
test_input[16496:16503] = '{32'hc188076f, 32'hc1e8ce95, 32'h424dd375, 32'h41e22f18, 32'h424ffb9e, 32'hc0f855b5, 32'hc1a00e03, 32'h41da85ac};
test_label[2062] = '{32'hc1a00e03};
test_output[2062] = '{32'h4290ec8d};
/*############ DEBUG ############
test_input[16496:16503] = '{-17.0036289086, -29.1008708921, 51.4564994611, 28.272995002, 51.9957203937, -7.76046227718, -20.0068411196, 27.315269148};
test_label[2062] = '{-20.0068411196};
test_output[2062] = '{72.4620111631};
############ END DEBUG ############*/
test_input[16504:16511] = '{32'hc25ebc07, 32'h42916ec5, 32'hc2168a95, 32'hc2960ca4, 32'hc24ab435, 32'h4236ce5a, 32'h4092d332, 32'h405c3ce6};
test_label[2063] = '{32'h4236ce5a};
test_output[2063] = '{32'h41d81e5f};
/*############ DEBUG ############
test_input[16504:16511] = '{-55.6836196438, 72.7163468465, -37.6353345784, -75.0246851119, -50.6759818054, 45.7015169683, 4.58828071926, 3.44121684503};
test_label[2063] = '{45.7015169683};
test_output[2063] = '{27.0148298783};
############ END DEBUG ############*/
test_input[16512:16519] = '{32'hc285a0f7, 32'hc2bbb174, 32'hc13c67bb, 32'hc09cb229, 32'h419c2460, 32'hc22c258e, 32'hc099b43a, 32'h428fab3b};
test_label[2064] = '{32'hc285a0f7};
test_output[2064] = '{32'h430aa619};
/*############ DEBUG ############
test_input[16512:16519] = '{-66.814384093, -93.8465866865, -11.7753243899, -4.89674812668, 19.5177619476, -43.0366763026, -4.80325054159, 71.8344373192};
test_label[2064] = '{-66.814384093};
test_output[2064] = '{138.648821412};
############ END DEBUG ############*/
test_input[16520:16527] = '{32'hc285fc31, 32'hc1ffe282, 32'hc2af4d60, 32'h41299083, 32'h3f4a20ba, 32'h41e00207, 32'h42ae810e, 32'h429e9dc9};
test_label[2065] = '{32'h41299083};
test_output[2065] = '{32'h42994f2c};
/*############ DEBUG ############
test_input[16520:16527] = '{-66.992560477, -31.9855994093, -87.6511226396, 10.5977814042, 0.789561852992, 28.0009893759, 87.25205916, 79.3081757126};
test_label[2065] = '{10.5977814042};
test_output[2065] = '{76.6546325188};
############ END DEBUG ############*/
test_input[16528:16535] = '{32'h421fbdb3, 32'hc1d0b4b3, 32'h4273c9a9, 32'h412a9fcd, 32'h41d502ee, 32'h420f0617, 32'h413cfee1, 32'h424be357};
test_label[2066] = '{32'hc1d0b4b3};
test_output[2066] = '{32'h42ae1207};
/*############ DEBUG ############
test_input[16528:16535] = '{39.9352537234, -26.088232272, 60.9469321354, 10.6640138085, 26.6264313268, 35.7559477826, 11.812226356, 50.9720097591};
test_label[2066] = '{-26.088232272};
test_output[2066] = '{87.0352109599};
############ END DEBUG ############*/
test_input[16536:16543] = '{32'h420541af, 32'h42396139, 32'h4261df1b, 32'h428942bd, 32'h41d278bb, 32'h408706d9, 32'h42a5c1cf, 32'h42bed0d2};
test_label[2067] = '{32'h42396139};
test_output[2067] = '{32'h4244406b};
/*############ DEBUG ############
test_input[16536:16543] = '{33.3141434462, 46.3449454444, 56.4678748923, 68.6303487229, 26.3089509986, 4.21958600892, 82.8785331279, 95.4078487244};
test_label[2067] = '{46.3449454444};
test_output[2067] = '{49.0629068991};
############ END DEBUG ############*/
test_input[16544:16551] = '{32'hc22fd244, 32'hc2a9daaa, 32'h41cec111, 32'hc20fb06c, 32'h42c3a7ec, 32'h418aa089, 32'h42c1d230, 32'hc2948abf};
test_label[2068] = '{32'h418aa089};
test_output[2068] = '{32'h42a1abe5};
/*############ DEBUG ############
test_input[16544:16551] = '{-43.9553393521, -84.9270803648, 25.844270677, -35.9222878816, 97.8279737505, 17.3283862965, 96.9105213714, -74.2709866641};
test_label[2068] = '{17.3283862965};
test_output[2068] = '{80.8357279292};
############ END DEBUG ############*/
test_input[16552:16559] = '{32'hc271bb4c, 32'h40bbfe73, 32'h428ea38e, 32'h42c3f96b, 32'h427c1dd5, 32'h420e76d2, 32'h429742c7, 32'hc2863f08};
test_label[2069] = '{32'hc271bb4c};
test_output[2069] = '{32'h431e6b89};
/*############ DEBUG ############
test_input[16552:16559] = '{-60.4329084781, 5.8748106013, 71.3194438729, 97.9871438156, 63.0291320712, 35.6160359716, 75.6304231281, -67.123111694};
test_label[2069] = '{-60.4329084781};
test_output[2069] = '{158.420052294};
############ END DEBUG ############*/
test_input[16560:16567] = '{32'hc296e205, 32'h429c68d3, 32'h41b15414, 32'hc1b614af, 32'hc1f0d574, 32'hc230ca58, 32'hc2103d07, 32'h42060d0e};
test_label[2070] = '{32'hc1b614af};
test_output[2070] = '{32'h42c9edff};
/*############ DEBUG ############
test_input[16560:16567] = '{-75.4414424184, 78.2047351663, 22.1660533667, -22.760099975, -30.1042260752, -44.1975998172, -36.0595980808, 33.5127488327};
test_label[2070] = '{-22.760099975};
test_output[2070] = '{100.964835141};
############ END DEBUG ############*/
test_input[16568:16575] = '{32'h422b58eb, 32'hc29de11d, 32'hc249e34f, 32'h42123c46, 32'hc288ebbe, 32'hc2c49d97, 32'h4284a3a1, 32'h40268ab0};
test_label[2071] = '{32'h422b58eb};
test_output[2071] = '{32'h41bbdcac};
/*############ DEBUG ############
test_input[16568:16575] = '{42.8368342931, -78.9396774348, -50.4719810899, 36.5588606534, -68.4604377342, -98.3077901328, 66.319584117, 2.60221486351};
test_label[2071] = '{42.8368342931};
test_output[2071] = '{23.482749824};
############ END DEBUG ############*/
test_input[16576:16583] = '{32'h423bb0c6, 32'hc25bf52c, 32'hc20dedb1, 32'hc02aa2eb, 32'hc0d150b6, 32'h415cc275, 32'h42693a0b, 32'h428ae512};
test_label[2072] = '{32'hc0d150b6};
test_output[2072] = '{32'h4297fa20};
/*############ DEBUG ############
test_input[16576:16583] = '{46.9226297649, -54.9894264833, -35.4821220997, -2.6661938027, -6.54110235183, 13.7974750504, 58.3066809043, 69.4474065388};
test_label[2072] = '{-6.54110235183};
test_output[2072] = '{75.9885233999};
############ END DEBUG ############*/
test_input[16584:16591] = '{32'h41d733dc, 32'hc22eb8a4, 32'h42884130, 32'hc2a045f0, 32'hc269221a, 32'hc2b90df5, 32'hc0b843d1, 32'h42579669};
test_label[2073] = '{32'hc2a045f0};
test_output[2073] = '{32'h43144390};
/*############ DEBUG ############
test_input[16584:16591] = '{26.9003216603, -43.6803143362, 68.1273201815, -80.1365993058, -58.2833018073, -92.5272584716, -5.75827850953, 53.896886105};
test_label[2073] = '{-80.1365993058};
test_output[2073] = '{148.263920148};
############ END DEBUG ############*/
test_input[16592:16599] = '{32'hc2b932ee, 32'hc1f25434, 32'h42900d06, 32'h428a904e, 32'h41dc3c05, 32'hc288798a, 32'h42c5c5f8, 32'hbfc867dd};
test_label[2074] = '{32'h42900d06};
test_output[2074] = '{32'h41d6e3c5};
/*############ DEBUG ############
test_input[16592:16599] = '{-92.5994745853, -30.2911149363, 72.025439417, 69.2818482174, 27.5293071595, -68.2373788197, 98.8866558556, -1.56566967055};
test_label[2074] = '{72.025439417};
test_output[2074] = '{26.8612164387};
############ END DEBUG ############*/
test_input[16600:16607] = '{32'h4254acfc, 32'hc0aa989f, 32'hc22ca75f, 32'h42a77e00, 32'hc1d694b3, 32'h42604757, 32'hc2928ef1, 32'hc2ac8f37};
test_label[2075] = '{32'hc0aa989f};
test_output[2075] = '{32'h42b2278a};
/*############ DEBUG ############
test_input[16600:16607] = '{53.1689285135, -5.3311302926, -43.1634498678, 83.7460921891, -26.8226079695, 56.0696684357, -73.2791814951, -86.2797150623};
test_label[2075] = '{-5.3311302926};
test_output[2075] = '{89.0772224817};
############ END DEBUG ############*/
test_input[16608:16615] = '{32'hc114c6a1, 32'h41bc6d5f, 32'h417e69f1, 32'hc22acc6b, 32'h42753dbe, 32'hc28aa3f7, 32'h3f42fe89, 32'h4299c9bf};
test_label[2076] = '{32'hc28aa3f7};
test_output[2076] = '{32'h431236db};
/*############ DEBUG ############
test_input[16608:16615] = '{-9.2984935408, 23.553403942, 15.9008649539, -42.6996262168, 61.3102932527, -69.3202462604, 0.76169642571, 76.8940377734};
test_label[2076] = '{-69.3202462604};
test_output[2076] = '{146.214284204};
############ END DEBUG ############*/
test_input[16616:16623] = '{32'hc28a21c8, 32'h3eb08c1b, 32'h42acfb0f, 32'h42c0beb1, 32'hc2a36809, 32'hc28b3d8e, 32'h427dd344, 32'hc193b4b4};
test_label[2077] = '{32'hc193b4b4};
test_output[2077] = '{32'h42e5abe4};
/*############ DEBUG ############
test_input[16616:16623] = '{-69.0659800958, 0.344818928514, 86.490352242, 96.3724421997, -81.7031937829, -69.6202250155, 63.4563129676, -18.4632339723};
test_label[2077] = '{-18.4632339723};
test_output[2077] = '{114.835727252};
############ END DEBUG ############*/
test_input[16624:16631] = '{32'hc28fadc7, 32'hc09b2ec1, 32'h42932a33, 32'hc29d2c00, 32'hc287defc, 32'h415bee3f, 32'hc1bebcad, 32'hc2bfe728};
test_label[2078] = '{32'hc29d2c00};
test_output[2078] = '{32'h43182b1a};
/*############ DEBUG ############
test_input[16624:16631] = '{-71.8394066941, -4.84945706006, 73.5824240933, -78.5859341241, -67.9355166026, 13.7456653074, -23.8421260843, -95.9514744269};
test_label[2078] = '{-78.5859341241};
test_output[2078] = '{152.168358217};
############ END DEBUG ############*/
test_input[16632:16639] = '{32'hc19355d1, 32'h42999b91, 32'hc20ee897, 32'hc2bc9392, 32'h42c28cbc, 32'hc2063ec4, 32'h42655b0f, 32'h4057ad18};
test_label[2079] = '{32'h42c28cbc};
test_output[2079] = '{32'h30b0de87};
/*############ DEBUG ############
test_input[16632:16639] = '{-18.4169019713, 76.8038402144, -35.7271395485, -94.2882226276, 97.2748751908, -33.5612961151, 57.3389244845, 3.36993987507};
test_label[2079] = '{97.2748751908};
test_output[2079] = '{1.28689314843e-09};
############ END DEBUG ############*/
test_input[16640:16647] = '{32'hc13fac40, 32'h3f081483, 32'hc21f2d02, 32'hc261648b, 32'h41830124, 32'h4282124a, 32'hc28b4102, 32'h41af9253};
test_label[2080] = '{32'h4282124a};
test_output[2080] = '{32'h80000000};
/*############ DEBUG ############
test_input[16640:16647] = '{-11.9795529939, 0.531563012102, -39.7939519271, -56.3481871212, 16.3755569996, 65.0357175416, -69.6269699739, 21.9464467616};
test_label[2080] = '{65.0357175416};
test_output[2080] = '{-0.0};
############ END DEBUG ############*/
test_input[16648:16655] = '{32'hc186db73, 32'h422910fc, 32'hc131f564, 32'hc1b61946, 32'h41823492, 32'hc19a64bb, 32'hc2c3b020, 32'hc19e46bc};
test_label[2081] = '{32'h422910fc};
test_output[2081] = '{32'h2cb56600};
/*############ DEBUG ############
test_input[16648:16655] = '{-16.8571530382, 42.2665853515, -11.1224096635, -22.7623399275, 16.2756699485, -19.2991847731, -97.8439949178, -19.7845390819};
test_label[2081] = '{42.2665853515};
test_output[2081] = '{5.15565368177e-12};
############ END DEBUG ############*/
test_input[16656:16663] = '{32'hc219a5be, 32'h427adebf, 32'hc1c7ec19, 32'hc2c41d8b, 32'h429a5649, 32'hc0eb902c, 32'hc2097e04, 32'h42943455};
test_label[2082] = '{32'hc2c41d8b};
test_output[2082] = '{32'h432f4593};
/*############ DEBUG ############
test_input[16656:16663] = '{-38.4118595052, 62.7175253405, -24.9902823064, -98.0576990344, 77.1685293016, -7.361349291, -34.3730626134, 74.1022073115};
test_label[2082] = '{-98.0576990344};
test_output[2082] = '{175.271768211};
############ END DEBUG ############*/
test_input[16664:16671] = '{32'hc277a9ff, 32'hc28b6c7a, 32'hc24821a2, 32'h420903c1, 32'hc1a5b309, 32'h40c83563, 32'hc2223a68, 32'hc26b08a5};
test_label[2083] = '{32'hc2223a68};
test_output[2083] = '{32'h42959f14};
/*############ DEBUG ############
test_input[16664:16671] = '{-61.9160126778, -69.7118700562, -50.0328464078, 34.2536650148, -20.7124204377, 6.2565167454, -40.5570356005, -58.7584435178};
test_label[2083] = '{-40.5570356005};
test_output[2083] = '{74.8107006153};
############ END DEBUG ############*/
test_input[16672:16679] = '{32'hc1df9032, 32'hc22741ad, 32'h41a56f33, 32'h42bbc28b, 32'h4224c39c, 32'h42bfc703, 32'hc25155d7, 32'hc29264f4};
test_label[2084] = '{32'h42bbc28b};
test_output[2084] = '{32'h40089d9c};
/*############ DEBUG ############
test_input[16672:16679] = '{-27.9454084936, -41.814135392, 20.6792969072, 93.8799662971, 41.1910241189, 95.8886944072, -52.3338289281, -73.1971756129};
test_label[2084] = '{93.8799662971};
test_output[2084] = '{2.13461969528};
############ END DEBUG ############*/
test_input[16680:16687] = '{32'hc284c0ac, 32'hc2a2fce1, 32'h413f93b2, 32'h4162fe66, 32'h42b2caad, 32'h428c3fa9, 32'hc1a87ab8, 32'hc20fa393};
test_label[2085] = '{32'h428c3fa9};
test_output[2085] = '{32'h419a2c0f};
/*############ DEBUG ############
test_input[16680:16687] = '{-66.3763108327, -81.4939067101, 11.9735584924, 14.187108699, 89.3958527726, 70.1243394447, -21.0599215419, -35.9097394222};
test_label[2085] = '{70.1243394447};
test_output[2085] = '{19.2715133321};
############ END DEBUG ############*/
test_input[16688:16695] = '{32'h426c839a, 32'h42ac7680, 32'hc2134bc4, 32'h41f109f3, 32'hc234d391, 32'h418c2b78, 32'hc26faa8c, 32'h428b9af0};
test_label[2086] = '{32'h418c2b78};
test_output[2086] = '{32'h42896ba2};
/*############ DEBUG ############
test_input[16688:16695] = '{59.1285186088, 86.2314438325, -36.8239907286, 30.1298587138, -45.2066084456, 17.5212246836, -59.9165515442, 69.8026143109};
test_label[2086] = '{17.5212246836};
test_output[2086] = '{68.7102192222};
############ END DEBUG ############*/
test_input[16696:16703] = '{32'h4187ffb8, 32'h42c07554, 32'hc2bfed00, 32'hc265d28d, 32'h41a4341d, 32'hc2817587, 32'h405432f2, 32'h41cf5290};
test_label[2087] = '{32'hc2bfed00};
test_output[2087] = '{32'h4340312a};
/*############ DEBUG ############
test_input[16696:16703] = '{16.9998629152, 96.2291553205, -95.9628906506, -57.4556175689, 20.5254464061, -64.7295418032, 3.31560936473, 25.9153141666};
test_label[2087] = '{-95.9628906506};
test_output[2087] = '{192.192045971};
############ END DEBUG ############*/
test_input[16704:16711] = '{32'h42be5f46, 32'hc20dc886, 32'h3f23c6a5, 32'h419bd1f6, 32'hc28cc2aa, 32'h40db38d8, 32'hc23cc235, 32'h41e7b262};
test_label[2088] = '{32'h3f23c6a5};
test_output[2088] = '{32'h42bd17b9};
/*############ DEBUG ############
test_input[16704:16711] = '{95.1860823462, -35.4458254899, 0.639749809439, 19.4775195717, -70.3802051327, 6.85068871024, -47.1896563263, 28.9621005865};
test_label[2088] = '{0.639749809439};
test_output[2088] = '{94.5463325367};
############ END DEBUG ############*/
test_input[16712:16719] = '{32'h429a6f0e, 32'hc0b9328e, 32'hc1e29936, 32'hc29a60a6, 32'h426102a5, 32'h3fae64e3, 32'h42b40430, 32'hc1c82c32};
test_label[2089] = '{32'h426102a5};
test_output[2089] = '{32'h420705ba};
/*############ DEBUG ############
test_input[16712:16719] = '{77.2169032413, -5.787421426, -28.3248109363, -77.1887699285, 56.2525838876, 1.36245385723, 90.0081750975, -25.0215795688};
test_label[2089] = '{56.2525838876};
test_output[2089] = '{33.7555939948};
############ END DEBUG ############*/
test_input[16720:16727] = '{32'hc1e116c1, 32'hc296fe93, 32'hc0dd02c3, 32'hc0a3d3f2, 32'hc22c95c4, 32'h429213a0, 32'h42955e61, 32'hc1b8cf89};
test_label[2090] = '{32'hc22c95c4};
test_output[2090] = '{32'h42ec0389};
/*############ DEBUG ############
test_input[16720:16727] = '{-28.1361105945, -75.4972162264, -6.9065873281, -5.11962237896, -43.1462537187, 73.0383292391, 74.6843311148, -23.1013354372};
test_label[2090] = '{-43.1462537187};
test_output[2090] = '{118.006904486};
############ END DEBUG ############*/
test_input[16728:16735] = '{32'hc1afd798, 32'h418ae7b8, 32'h41c2957f, 32'hc2c5bff4, 32'h4244d3f1, 32'h41730f41, 32'hc225a46b, 32'h408c5d9f};
test_label[2091] = '{32'h408c5d9f};
test_output[2091] = '{32'h4233483d};
/*############ DEBUG ############
test_input[16728:16735] = '{-21.9802712357, 17.36314341, 24.3229969747, -98.874910848, 49.2069730187, 15.1912239827, -41.4105647809, 4.38642821557};
test_label[2091] = '{4.38642821557};
test_output[2091] = '{44.8205448032};
############ END DEBUG ############*/
test_input[16736:16743] = '{32'h4123bf90, 32'hc1cc01cd, 32'h42011fcc, 32'hc28a1d60, 32'hc10fb9bf, 32'hc2450bfe, 32'hc245120c, 32'hc14f9eb0};
test_label[2092] = '{32'hc1cc01cd};
test_output[2092] = '{32'h426720b3};
/*############ DEBUG ############
test_input[16736:16743] = '{10.2342677911, -25.5008798727, 32.2810514877, -69.0573759429, -8.98284774832, -49.2617105472, -49.2676257399, -12.9762421316};
test_label[2092] = '{-25.5008798727};
test_output[2092] = '{57.7819313607};
############ END DEBUG ############*/
test_input[16744:16751] = '{32'h42921554, 32'h4155422f, 32'h42c4c346, 32'hc2311bac, 32'h41c0d0bc, 32'h4107ce94, 32'hc10a2750, 32'h42b9aab3};
test_label[2093] = '{32'h42921554};
test_output[2093] = '{32'h41cabfbf};
/*############ DEBUG ############
test_input[16744:16751] = '{73.0416574173, 13.3286579806, 98.3813955524, -44.2770236897, 24.1019215972, 8.48793386614, -8.63459802409, 92.8333994923};
test_label[2093] = '{73.0416574173};
test_output[2093] = '{25.3436258235};
############ END DEBUG ############*/
test_input[16752:16759] = '{32'hc18f9128, 32'hc1f2e97e, 32'h42af0318, 32'h41f06149, 32'h4275a155, 32'h401e7c71, 32'hc112599a, 32'hc283475e};
test_label[2094] = '{32'hc283475e};
test_output[2094] = '{32'h4319253b};
/*############ DEBUG ############
test_input[16752:16759] = '{-17.9458774416, -30.3640092179, 87.5060428023, 30.0475023862, 61.4075501188, 2.47634536849, -9.14687540448, -65.6393924409};
test_label[2094] = '{-65.6393924409};
test_output[2094] = '{153.145435243};
############ END DEBUG ############*/
test_input[16760:16767] = '{32'h42313aca, 32'h42be6a7a, 32'hc25dfac9, 32'hc20eed5c, 32'hc24f3fc2, 32'hbeb6adb5, 32'hc1025dee, 32'h427ba894};
test_label[2095] = '{32'h427ba894};
test_output[2095] = '{32'h42012c61};
/*############ DEBUG ############
test_input[16760:16767] = '{44.3074107328, 95.2079652704, -55.4949074824, -35.7317959582, -51.8122632542, -0.356794039825, -8.14793228669, 62.9146280719};
test_label[2095] = '{62.9146280719};
test_output[2095] = '{32.2933371985};
############ END DEBUG ############*/
test_input[16768:16775] = '{32'hc0b461c6, 32'hc24a89fa, 32'h410503b6, 32'h4203a1e4, 32'h423f969b, 32'h42a8f55e, 32'h428b4797, 32'hc2c5f365};
test_label[2096] = '{32'h428b4797};
test_output[2096] = '{32'h416d6e35};
/*############ DEBUG ############
test_input[16768:16775] = '{-5.63693521159, -50.6347440733, 8.3134055933, 32.9080954842, 47.897075199, 84.4792331541, 69.6398275273, -98.9753808227};
test_label[2096] = '{69.6398275273};
test_output[2096] = '{14.839405986};
############ END DEBUG ############*/
test_input[16776:16783] = '{32'h41a9923d, 32'hc2920eae, 32'h42577b63, 32'h41e8e5e2, 32'hc20465ee, 32'h41cb2f82, 32'hc2c14aa9, 32'hc2b68c9d};
test_label[2097] = '{32'h42577b63};
test_output[2097] = '{32'h2d9f6b00};
/*############ DEBUG ############
test_input[16776:16783] = '{21.1964055897, -73.0286726245, 53.8704953857, 29.1122483065, -33.0995411833, 25.3981967659, -96.6458216931, -91.274638759};
test_label[2097] = '{53.8704953857};
test_output[2097] = '{1.81237247434e-11};
############ END DEBUG ############*/
test_input[16784:16791] = '{32'hc2750cdc, 32'h422ae1f3, 32'h42261996, 32'h428a9ff0, 32'hc28fd44b, 32'h41b29454, 32'hc28f24ef, 32'hc2c5ca92};
test_label[2098] = '{32'hc2750cdc};
test_output[2098] = '{32'h4302932f};
/*############ DEBUG ############
test_input[16784:16791] = '{-61.2625575048, 42.7206537877, 41.5249853213, 69.3123741298, -71.9146336049, 22.3224254054, -71.5721385453, -98.8956449998};
test_label[2098] = '{-61.2625575048};
test_output[2098] = '{130.574931635};
############ END DEBUG ############*/
test_input[16792:16799] = '{32'hc19eb82a, 32'h41e461b0, 32'hc1d3b900, 32'hc259c75f, 32'hc1cb971b, 32'hc1929a3b, 32'hc0313355, 32'h420ec3ef};
test_label[2099] = '{32'h420ec3ef};
test_output[2099] = '{32'h3a4efa4c};
/*############ DEBUG ############
test_input[16792:16799] = '{-19.839923555, 28.5476993044, -26.4653311676, -54.444699663, -25.4487814284, -18.325306978, -2.76875796292, 35.6913425799};
test_label[2099] = '{35.6913425799};
test_output[2099] = '{0.000789557354652};
############ END DEBUG ############*/
test_input[16800:16807] = '{32'h413e5072, 32'h425f2fca, 32'hc28457f2, 32'hc1cc2ebe, 32'h42c7308f, 32'h42a0f1d7, 32'h4099bda1, 32'h42567ea7};
test_label[2100] = '{32'h42567ea7};
test_output[2100] = '{32'h4237e276};
/*############ DEBUG ############
test_input[16800:16807] = '{11.894640398, 55.7966683998, -66.171767986, -25.5228228984, 99.5948375894, 80.4723425014, 4.80439821047, 53.6236839346};
test_label[2100] = '{53.6236839346};
test_output[2100] = '{45.9711536597};
############ END DEBUG ############*/
test_input[16808:16815] = '{32'hc28ff0d1, 32'hbd937bd3, 32'hc2b5f1c8, 32'h4290e825, 32'hc1a09383, 32'h42bae213, 32'hc1a27d02, 32'h41b907a0};
test_label[2101] = '{32'hc28ff0d1};
test_output[2101] = '{32'h43256972};
/*############ DEBUG ############
test_input[16808:16815] = '{-71.9703421864, -0.0720135188198, -90.9722263618, 72.4534055135, -20.072027158, 93.441548355, -20.3110393388, 23.1287234314};
test_label[2101] = '{-71.9703421864};
test_output[2101] = '{165.411890542};
############ END DEBUG ############*/
test_input[16816:16823] = '{32'hc2c70265, 32'hc1a151dc, 32'hc20a6296, 32'hc2a4c1f7, 32'h41b253d6, 32'h428b1445, 32'h413bee3a, 32'hbf632625};
test_label[2102] = '{32'hc1a151dc};
test_output[2102] = '{32'h42b368bc};
/*############ DEBUG ############
test_input[16816:16823] = '{-99.5046742995, -20.164970499, -34.596275938, -82.3788378529, 22.2909348999, 69.5395857981, 11.7456608868, -0.88730079779};
test_label[2102] = '{-20.164970499};
test_output[2102] = '{89.7045562971};
############ END DEBUG ############*/
test_input[16824:16831] = '{32'hc25a7723, 32'h41c9ea1f, 32'h41c091b2, 32'h426ca606, 32'h425a6a61, 32'hc11c6ebc, 32'h420bad36, 32'h4210bc82};
test_label[2103] = '{32'h426ca606};
test_output[2103] = '{32'h3c2ad148};
/*############ DEBUG ############
test_input[16824:16831] = '{-54.6163443039, 25.2393174757, 24.0711402335, 59.1621333063, 54.60388597, -9.77703440334, 34.9191511398, 36.1840880628};
test_label[2103] = '{59.1621333063};
test_output[2103] = '{0.0104258728412};
############ END DEBUG ############*/
test_input[16832:16839] = '{32'h42b2cd66, 32'hc1f70a56, 32'h42a68ff9, 32'hc2a6b4d9, 32'hc27752eb, 32'h41dbbfd5, 32'h4294026d, 32'hc2aae9c1};
test_label[2104] = '{32'hc2a6b4d9};
test_output[2104] = '{32'h432cc1b0};
/*############ DEBUG ############
test_input[16832:16839] = '{89.4011713505, -30.8800462073, 83.2811981643, -83.3532167876, -61.8309730349, 27.4686675553, 74.0047351138, -85.456552254};
test_label[2104] = '{-83.3532167876};
test_output[2104] = '{172.756584445};
############ END DEBUG ############*/
test_input[16840:16847] = '{32'h42711fe5, 32'hc22d3d08, 32'h41873193, 32'h4292e0eb, 32'hc2c5253d, 32'h42226ba9, 32'hc2283bde, 32'h4210aa91};
test_label[2105] = '{32'h42711fe5};
test_output[2105] = '{32'h415287c2};
/*############ DEBUG ############
test_input[16840:16847] = '{60.281147577, -43.3096027345, 16.8992059231, 73.4392895198, -98.5727298451, 40.6051351334, -42.0584628952, 36.1665706535};
test_label[2105] = '{60.281147577};
test_output[2105] = '{13.1581438726};
############ END DEBUG ############*/
test_input[16848:16855] = '{32'h427eb269, 32'hc15843a7, 32'hc2959403, 32'h42571de0, 32'hc24218d8, 32'hc2bec7b7, 32'hc259f9cc, 32'h42254292};
test_label[2106] = '{32'h427eb269};
test_output[2106] = '{32'h38537ca3};
/*############ DEBUG ############
test_input[16848:16855] = '{63.6742281722, -13.5165162813, -74.7890825958, 53.7791744605, -48.5242633187, -95.390067811, -54.493941156, 41.3150094059};
test_label[2106] = '{63.6742281722};
test_output[2106] = '{5.04223988259e-05};
############ END DEBUG ############*/
test_input[16856:16863] = '{32'h41c686de, 32'hc2c4550e, 32'hc0863be0, 32'hc2af7b1b, 32'hc2421686, 32'h423b5df3, 32'h4107e600, 32'hc2560ac6};
test_label[2107] = '{32'hc0863be0};
test_output[2107] = '{32'h424c256f};
/*############ DEBUG ############
test_input[16856:16863] = '{24.8158527007, -98.166124568, -4.19480894226, -87.7404431481, -48.5219963715, 46.8417463429, 8.49365213933, -53.510521352};
test_label[2107] = '{-4.19480894226};
test_output[2107] = '{51.0365552854};
############ END DEBUG ############*/
test_input[16864:16871] = '{32'h411cd50a, 32'hc2b602e5, 32'hc2aa3985, 32'hc20bb164, 32'h424425c1, 32'hc2959a4f, 32'h421bd61c, 32'hbc852781};
test_label[2108] = '{32'hc20bb164};
test_output[2108] = '{32'h42a7eb98};
/*############ DEBUG ############
test_input[16864:16871] = '{9.80201141007, -91.0056518128, -85.1123427886, -34.9232340315, 49.0368695362, -74.8013848665, 38.9590928445, -0.0162541886739};
test_label[2108] = '{-34.9232340315};
test_output[2108] = '{83.9601455695};
############ END DEBUG ############*/
test_input[16872:16879] = '{32'hc228d77d, 32'hc1cae32c, 32'h4277e259, 32'h425dd09e, 32'hc29193e7, 32'hc2584540, 32'h42aba2f4, 32'hc2a844a8};
test_label[2109] = '{32'hc1cae32c};
test_output[2109] = '{32'h42de5bbf};
/*############ DEBUG ############
test_input[16872:16879] = '{-42.2104371949, -25.3609229243, 61.9710434647, 55.4537288965, -72.7888715344, -54.0676259219, 85.8182703143, -84.1340969562};
test_label[2109] = '{-25.3609229243};
test_output[2109] = '{111.179193239};
############ END DEBUG ############*/
test_input[16880:16887] = '{32'h42af52d1, 32'h42c1fe47, 32'h42a31147, 32'h42509af8, 32'h4191ae25, 32'hc2a3a757, 32'h42c1808b, 32'hc23ba897};
test_label[2110] = '{32'h42c1fe47};
test_output[2110] = '{32'h3f13f310};
/*############ DEBUG ############
test_input[16880:16887] = '{87.6617485263, 96.996636516, 81.5337458074, 52.1513378655, 18.2100312124, -81.8268351424, 96.751058719, -46.9146366737};
test_label[2110] = '{96.996636516};
test_output[2110] = '{0.577927616418};
############ END DEBUG ############*/
test_input[16888:16895] = '{32'hc2b64caa, 32'h418f9fe7, 32'hc23dd7b4, 32'h408628a6, 32'hc2ab3543, 32'hc157ecf9, 32'hc24e2514, 32'hc20bcace};
test_label[2111] = '{32'hc2b64caa};
test_output[2111] = '{32'h42da34a4};
/*############ DEBUG ############
test_input[16888:16895] = '{-91.1497382571, 17.9530765854, -47.4606462871, 4.19246196693, -85.6040271996, -13.4953541758, -51.5362089223, -34.9480517313};
test_label[2111] = '{-91.1497382571};
test_output[2111] = '{109.102815899};
############ END DEBUG ############*/
test_input[16896:16903] = '{32'hc2af3fad, 32'h42901f90, 32'h420a62bf, 32'hc2893fcf, 32'hc202733c, 32'h42bba4b3, 32'hc20f00a0, 32'hc1b345fc};
test_label[2112] = '{32'hc20f00a0};
test_output[2112] = '{32'h43019281};
/*############ DEBUG ############
test_input[16896:16903] = '{-87.6243689006, 72.0616422546, 34.5964332281, -68.6246226134, -32.6125337545, 93.8216767853, -35.7506096859, -22.409172992};
test_label[2112] = '{-35.7506096859};
test_output[2112] = '{129.572286472};
############ END DEBUG ############*/
test_input[16904:16911] = '{32'h4187066f, 32'hc2c3dbfb, 32'hc221c669, 32'h41dccd77, 32'h41984e40, 32'hc2c6dc77, 32'h4274dbdc, 32'h416a5f25};
test_label[2113] = '{32'hc2c3dbfb};
test_output[2113] = '{32'h431f24f4};
/*############ DEBUG ############
test_input[16904:16911] = '{16.878140599, -97.9296465123, -40.4437602778, 27.6003241992, 19.038208775, -99.430592448, 61.2147067664, 14.6482281998};
test_label[2113] = '{-97.9296465123};
test_output[2113] = '{159.144353279};
############ END DEBUG ############*/
test_input[16912:16919] = '{32'h423b02c8, 32'h41d71e94, 32'h42568406, 32'h42297909, 32'h411a01da, 32'h42826fef, 32'hc25e1d16, 32'h4199fe9f};
test_label[2114] = '{32'h42297909};
test_output[2114] = '{32'h41b6cdae};
/*############ DEBUG ############
test_input[16912:16919] = '{46.7527144768, 26.8899308168, 53.6289303105, 42.3681989419, 9.62545248608, 65.2186182548, -55.5284050767, 19.2493260248};
test_label[2114] = '{42.3681989419};
test_output[2114] = '{22.8504285836};
############ END DEBUG ############*/
test_input[16920:16927] = '{32'h42484287, 32'h4254450f, 32'h4273ce55, 32'hc2bbec94, 32'hc2ae4ecb, 32'hc2821c00, 32'hc2b3f34d, 32'hc2991a78};
test_label[2115] = '{32'h4254450f};
test_output[2115] = '{32'h40fc4d69};
/*############ DEBUG ############
test_input[16920:16927] = '{50.064968036, 53.0674416339, 60.9514956276, -93.9620632634, -87.1538944643, -65.0546869472, -89.9751996704, -76.5516939177};
test_label[2115] = '{53.0674416339};
test_output[2115] = '{7.88444932687};
############ END DEBUG ############*/
test_input[16928:16935] = '{32'hbf26e2f2, 32'h42bcd6e7, 32'hc2bbd780, 32'hc2868ff1, 32'hc20385b3, 32'h422b0cf0, 32'hc26ecf0b, 32'h42b87c49};
test_label[2116] = '{32'h42b87c49};
test_output[2116] = '{32'h40123377};
/*############ DEBUG ############
test_input[16928:16935] = '{-0.65190041988, 94.4197335918, -93.9209010886, -67.2811339566, -32.8805649872, 42.7626351989, -59.7021896051, 92.2427451565};
test_label[2116] = '{92.2427451565};
test_output[2116] = '{2.28439109249};
############ END DEBUG ############*/
test_input[16936:16943] = '{32'h426b89e2, 32'hc1bc2f6a, 32'h425e3cb3, 32'h423a44b5, 32'hc2637659, 32'hc11619b9, 32'hc2918af2, 32'h42964492};
test_label[2117] = '{32'hc2637659};
test_output[2117] = '{32'h4303ffdf};
/*############ DEBUG ############
test_input[16936:16943] = '{58.88464966, -23.5231516305, 55.559275811, 46.5670951194, -56.8655753192, -9.38128015343, -72.7713750318, 75.1339246309};
test_label[2117] = '{-56.8655753192};
test_output[2117] = '{131.999500041};
############ END DEBUG ############*/
test_input[16944:16951] = '{32'h42ad4575, 32'h410f41dd, 32'h42a617af, 32'hc12a8115, 32'h4292381e, 32'h418c74de, 32'h41868988, 32'hc20c3d8c};
test_label[2118] = '{32'h42ad4575};
test_output[2118] = '{32'h3cdf2a01};
/*############ DEBUG ############
test_input[16944:16951] = '{86.6356606259, 8.95357951807, 83.04625795, -10.6565143314, 73.109604859, 17.557063539, 16.8171541431, -35.0601027704};
test_label[2118] = '{86.6356606259};
test_output[2118] = '{0.0272417083885};
############ END DEBUG ############*/
test_input[16952:16959] = '{32'hc2275fb5, 32'h402acf2d, 32'h4231a743, 32'h42c687a3, 32'h42afad12, 32'hc20c9a7c, 32'h420a078a, 32'hc1a3cb80};
test_label[2119] = '{32'h420a078a};
test_output[2119] = '{32'h428183df};
/*############ DEBUG ############
test_input[16952:16959] = '{-41.8434637645, 2.66889501625, 44.4133421629, 99.2649120799, 87.8380281063, -35.1508651268, 34.5073627145, -20.4743649025};
test_label[2119] = '{34.5073627145};
test_output[2119] = '{64.7575602639};
############ END DEBUG ############*/
test_input[16960:16967] = '{32'h421a8951, 32'h410c936e, 32'h4156702b, 32'h41b46e07, 32'hbeb8fa53, 32'hc2c3176c, 32'hc210891a, 32'h42b18284};
test_label[2120] = '{32'h421a8951};
test_output[2120] = '{32'h42487bb7};
/*############ DEBUG ############
test_input[16960:16967] = '{38.6340971283, 8.78599371709, 13.4023847083, 22.5537240497, -0.361284822355, -97.5457453835, -36.13388893, 88.7549126165};
test_label[2120] = '{38.6340971283};
test_output[2120] = '{50.1208154882};
############ END DEBUG ############*/
test_input[16968:16975] = '{32'hc1a4e3c2, 32'hc206f489, 32'h428c195b, 32'hc18c9975, 32'hc2adb55c, 32'h41791440, 32'hc2395a48, 32'h4169ed0f};
test_label[2121] = '{32'hc2adb55c};
test_output[2121] = '{32'h431ce75b};
/*############ DEBUG ############
test_input[16968:16975] = '{-20.6112103302, -33.7388041723, 70.0495224044, -17.5749307506, -86.8542169217, 15.5674441625, -46.3381646171, 14.6203759476};
test_label[2121] = '{-86.8542169217};
test_output[2121] = '{156.903739326};
############ END DEBUG ############*/
test_input[16976:16983] = '{32'h423dbcbb, 32'h4286901b, 32'h42a51a1b, 32'hc1e6ed89, 32'hc130cd30, 32'hc20bdb02, 32'hc29920d9, 32'hc27ed4b4};
test_label[2122] = '{32'h423dbcbb};
test_output[2122] = '{32'h420c777c};
/*############ DEBUG ############
test_input[16976:16983] = '{47.4343061394, 67.2814567556, 82.5509883082, -28.8659846654, -11.0500946974, -34.9638766654, -76.564158952, -63.7077187097};
test_label[2122] = '{47.4343061394};
test_output[2122] = '{35.1166824024};
############ END DEBUG ############*/
test_input[16984:16991] = '{32'h40ea1ed0, 32'h422109ed, 32'h41b18077, 32'hc2183898, 32'h42126607, 32'h415e5830, 32'h42af83d2, 32'h425a51d2};
test_label[2123] = '{32'h415e5830};
test_output[2123] = '{32'h4293b8cc};
/*############ DEBUG ############
test_input[16984:16991] = '{7.31626131899, 40.2596913791, 22.1877266968, -38.0552658625, 36.5996361979, 13.8965303804, 87.7574644211, 54.5799017508};
test_label[2123] = '{13.8965303804};
test_output[2123] = '{73.8609340407};
############ END DEBUG ############*/
test_input[16992:16999] = '{32'h426cd8d2, 32'hc2917063, 32'hc20319d8, 32'hc2135f93, 32'h41ca4a6b, 32'hc279b7f1, 32'hc11e9ee0, 32'h41581456};
test_label[2124] = '{32'h41ca4a6b};
test_output[2124] = '{32'h4207b39d};
/*############ DEBUG ############
test_input[16992:16999] = '{59.2117394333, -72.7195045766, -32.7752398559, -36.8433343971, 25.2863373948, -62.4296308613, -9.91378831655, 13.5049646703};
test_label[2124] = '{25.2863373948};
test_output[2124] = '{33.9254020385};
############ END DEBUG ############*/
test_input[17000:17007] = '{32'hc273c051, 32'h42a6d5fc, 32'hc28b7551, 32'h3fa4435f, 32'h42a0c8de, 32'h420d7d16, 32'h41e443af, 32'h414f408e};
test_label[2125] = '{32'h41e443af};
test_output[2125] = '{32'h425bbaa7};
/*############ DEBUG ############
test_input[17000:17007] = '{-60.9378077679, 83.417939079, -69.729131246, 1.2833059668, 80.3923211977, 35.3721556847, 28.5330483156, 12.9532606085};
test_label[2125] = '{28.5330483156};
test_output[2125] = '{54.9322778748};
############ END DEBUG ############*/
test_input[17008:17015] = '{32'h41c1292a, 32'h420334f9, 32'hc2829988, 32'h42328b93, 32'h41ca722f, 32'h41570961, 32'hc290d726, 32'h424eff0f};
test_label[2126] = '{32'h424eff0f};
test_output[2126] = '{32'h3a5576f4};
/*############ DEBUG ############
test_input[17008:17015] = '{24.1451004804, 32.8017296689, -65.2998677923, 44.636302554, 25.3057530431, 13.4397896097, -72.4202101172, 51.7490806016};
test_label[2126] = '{51.7490806016};
test_output[2126] = '{0.00081430304349};
############ END DEBUG ############*/
test_input[17016:17023] = '{32'h42a5a2c6, 32'hc287344e, 32'hc2c0b0ec, 32'h41bc7d8f, 32'h4286e656, 32'h42b1eb5c, 32'h40eeb955, 32'h4116ed62};
test_label[2127] = '{32'h42a5a2c6};
test_output[2127] = '{32'h40c49af8};
/*############ DEBUG ############
test_input[17016:17023] = '{82.8179152618, -67.6021567028, -96.3455521076, 23.5613079414, 67.4498734947, 88.9596833888, 7.46012374479, 9.43295436431};
test_label[2127] = '{82.8179152618};
test_output[2127] = '{6.14391693394};
############ END DEBUG ############*/
test_input[17024:17031] = '{32'h414f9837, 32'h41b246e2, 32'hc197abc3, 32'hc1f8ce03, 32'h42c58594, 32'h42964438, 32'hc1d53188, 32'hc21f3eef};
test_label[2128] = '{32'h42964438};
test_output[2128] = '{32'h41bd0572};
/*############ DEBUG ############
test_input[17024:17031] = '{12.9746619951, 22.2846108082, -18.9588671252, -31.1005921728, 98.7608970262, 75.1332372805, -26.6491853228, -39.8114585207};
test_label[2128] = '{75.1332372805};
test_output[2128] = '{23.6276597457};
############ END DEBUG ############*/
test_input[17032:17039] = '{32'h4221ba68, 32'hc253407e, 32'hc2c0289e, 32'h418f5399, 32'hc2bd4599, 32'hc26ca6a1, 32'hc2be125c, 32'h412fb0f8};
test_label[2129] = '{32'h418f5399};
test_output[2129] = '{32'h41b42137};
/*############ DEBUG ############
test_input[17032:17039] = '{40.4320372662, -52.812982452, -96.0793294422, 17.915819282, -94.6359293113, -59.1627251713, -95.035861014, 10.9807056903};
test_label[2129] = '{17.915819282};
test_output[2129] = '{22.5162179843};
############ END DEBUG ############*/
test_input[17040:17047] = '{32'hc27a6eeb, 32'h41dc8f99, 32'h4210e098, 32'h420c3997, 32'h3ff2999d, 32'hc2ae6b46, 32'hc237fdbf, 32'hc270437e};
test_label[2130] = '{32'h4210e098};
test_output[2130] = '{32'h3e8b4e46};
/*############ DEBUG ############
test_input[17040:17047] = '{-62.6083168783, 27.5701155693, 36.2193293666, 35.0562386407, 1.89531291588, -87.2095210764, -45.9978002311, -60.0659112012};
test_label[2130] = '{36.2193293666};
test_output[2130] = '{0.272081545609};
############ END DEBUG ############*/
test_input[17048:17055] = '{32'h42b6ce51, 32'h418a725c, 32'hc290437e, 32'h42514a3a, 32'h42a3bc84, 32'hc14658c7, 32'hc2410961, 32'h4293039a};
test_label[2131] = '{32'hc290437e};
test_output[2131] = '{32'h432388ec};
/*############ DEBUG ############
test_input[17048:17055] = '{91.4029625769, 17.3058388221, -72.1318226762, 52.3224875324, 81.8681919885, -12.3966738107, -48.259160355, 73.5070316245};
test_label[2131] = '{-72.1318226762};
test_output[2131] = '{163.534857561};
############ END DEBUG ############*/
test_input[17056:17063] = '{32'h41e3a4fe, 32'h42aa736e, 32'hc2a9074e, 32'hc29b6ac0, 32'h3f36e198, 32'h42bbf9f4, 32'hc22ecef3, 32'hc2b62d02};
test_label[2132] = '{32'hc29b6ac0};
test_output[2132] = '{32'h432bb264};
/*############ DEBUG ############
test_input[17056:17063] = '{28.455562469, 85.2254453044, -84.5142688166, -77.7084930515, 0.714379767829, 93.9881874201, -43.7020994902, -91.0879092434};
test_label[2132] = '{-77.7084930515};
test_output[2132] = '{171.696836914};
############ END DEBUG ############*/
test_input[17064:17071] = '{32'hc25d0fd5, 32'h4211ab09, 32'hc286a9c6, 32'h42a09b28, 32'hc22bea7e, 32'hc2a900f4, 32'hc231239c, 32'hc18053eb};
test_label[2133] = '{32'hc231239c};
test_output[2133] = '{32'h42f92cf6};
/*############ DEBUG ############
test_input[17064:17071] = '{-55.2654611805, 36.417026828, -67.3315897626, 80.3030401389, -42.9789971498, -84.5018593333, -44.2847754736, -16.0409752138};
test_label[2133] = '{-44.2847754736};
test_output[2133] = '{124.587815612};
############ END DEBUG ############*/
test_input[17072:17079] = '{32'h42235958, 32'hc1ae7c1c, 32'h42307443, 32'hc21bf28c, 32'hc262c4f4, 32'hbf290f3a, 32'h4259ab2f, 32'hc28fe18b};
test_label[2134] = '{32'hc262c4f4};
test_output[2134] = '{32'h42de3816};
/*############ DEBUG ############
test_input[17072:17079] = '{40.8372514545, -21.8106010082, 44.1135373514, -38.9868603727, -56.6923367138, -0.660388603649, 54.4171706647, -71.9405149174};
test_label[2134] = '{-56.6923367138};
test_output[2134] = '{111.109542155};
############ END DEBUG ############*/
test_input[17080:17087] = '{32'hc226a84e, 32'hc18efba9, 32'hc223b16a, 32'hc27b9d19, 32'hc2ae2676, 32'hc2a81268, 32'hc24baa8c, 32'h41e62fc4};
test_label[2135] = '{32'hc18efba9};
test_output[2135] = '{32'h423a95b7};
/*############ DEBUG ############
test_input[17080:17087] = '{-41.6643599639, -17.8728815898, -40.9232553752, -62.9034170355, -87.0751210152, -84.035948652, -50.9165492703, 28.7733229769};
test_label[2135] = '{-17.8728815898};
test_output[2135] = '{46.6462045667};
############ END DEBUG ############*/
test_input[17088:17095] = '{32'h429a2694, 32'h3f99abe4, 32'h4226ffcf, 32'hbfb40496, 32'h41222fdc, 32'hc2c6a36b, 32'hc2884f98, 32'hc29ee451};
test_label[2136] = '{32'hc2884f98};
test_output[2136] = '{32'h43113b16};
/*############ DEBUG ############
test_input[17088:17095] = '{77.0753491252, 1.20055820159, 41.7498138152, -1.40638992735, 10.1366845875, -99.3191775658, -68.1554586072, -79.4459285154};
test_label[2136] = '{-68.1554586072};
test_output[2136] = '{145.230807732};
############ END DEBUG ############*/
test_input[17096:17103] = '{32'h42157f78, 32'hc10ea164, 32'h42a770c5, 32'h429faf6e, 32'h42a16e21, 32'hc2b767c9, 32'h42c3b830, 32'h422f1d78};
test_label[2137] = '{32'h429faf6e};
test_output[2137] = '{32'h4190230b};
/*############ DEBUG ############
test_input[17096:17103] = '{37.3744807457, -8.91440206204, 83.7202522253, 79.8426331756, 80.7150953986, -91.7027073567, 97.8597435635, 43.7787775403};
test_label[2137] = '{79.8426331756};
test_output[2137] = '{18.017111162};
############ END DEBUG ############*/
test_input[17104:17111] = '{32'hc2ab5b7c, 32'hc2609859, 32'h418420bd, 32'h402b58a8, 32'hc27a82b6, 32'hc26d0d55, 32'hc26d3830, 32'hc22b5439};
test_label[2138] = '{32'hc2609859};
test_output[2138] = '{32'h4291545c};
/*############ DEBUG ############
test_input[17104:17111] = '{-85.6786833056, -56.1487783362, 16.5159859305, 2.67728611666, -62.6276474278, -59.2630210101, -59.3048692739, -42.8322503953};
test_label[2138] = '{-56.1487783362};
test_output[2138] = '{72.6647652437};
############ END DEBUG ############*/
test_input[17112:17119] = '{32'h429d2653, 32'hc23cb64a, 32'h424d1b7c, 32'h42057ffb, 32'h4253dcdd, 32'h42a7928d, 32'h42b7f339, 32'h4277f751};
test_label[2139] = '{32'hc23cb64a};
test_output[2139] = '{32'h430b2741};
/*############ DEBUG ############
test_input[17112:17119] = '{78.5748554356, -47.1780158352, 51.2768416537, 33.3749813013, 52.9656886649, 83.7862297469, 91.9750415806, 61.9915202713};
test_label[2139] = '{-47.1780158352};
test_output[2139] = '{139.153336635};
############ END DEBUG ############*/
test_input[17120:17127] = '{32'h411b34e6, 32'h4076ac92, 32'h4294b868, 32'hc2842e5f, 32'hc2a95e6a, 32'hc174c824, 32'hc1a80067, 32'hc2a92937};
test_label[2140] = '{32'h4294b868};
test_output[2140] = '{32'h80000000};
/*############ DEBUG ############
test_input[17120:17127] = '{9.70041496327, 3.85428285423, 74.3601685659, -66.0905649948, -84.6844034545, -15.2988625297, -21.0001970277, -84.5804961618};
test_label[2140] = '{74.3601685659};
test_output[2140] = '{-0.0};
############ END DEBUG ############*/
test_input[17128:17135] = '{32'hc2c42ce6, 32'h42afa852, 32'hc0816af9, 32'hc27476f1, 32'hc1e1190c, 32'hc28f18e5, 32'h4250c01b, 32'h427ad591};
test_label[2141] = '{32'hc2c42ce6};
test_output[2141] = '{32'h4339ea9c};
/*############ DEBUG ############
test_input[17128:17135] = '{-98.0876933912, 87.8287518313, -4.04430805906, -61.1161519292, -28.1372296903, -71.5486219333, 52.1876022789, 62.7085614887};
test_label[2141] = '{-98.0876933912};
test_output[2141] = '{185.916445223};
############ END DEBUG ############*/
test_input[17136:17143] = '{32'hc200d728, 32'h429507db, 32'h3fe7b414, 32'hc299e998, 32'h42526aa7, 32'hc29995c3, 32'h422ceeb7, 32'hc287fe57};
test_label[2142] = '{32'hc287fe57};
test_output[2142] = '{32'h430e8319};
/*############ DEBUG ############
test_input[17136:17143] = '{-32.2101142894, 74.5153453706, 1.81018304551, -76.9562384918, 52.6041540615, -76.792503624, 43.2331187615, -67.9967548454};
test_label[2142] = '{-67.9967548454};
test_output[2142] = '{142.512100216};
############ END DEBUG ############*/
test_input[17144:17151] = '{32'hc223c295, 32'h40899aed, 32'hc2c64c11, 32'hc29e6fa3, 32'h42368a1a, 32'hc2b17bbe, 32'h428b1240, 32'h41e68363};
test_label[2143] = '{32'h41e68363};
test_output[2143] = '{32'h4222e2ce};
/*############ DEBUG ############
test_input[17144:17151] = '{-40.9400225524, 4.30016197188, -99.1485637367, -79.2180377105, 45.6348653902, -88.7416872209, 69.5356444227, 28.8141540879};
test_label[2143] = '{28.8141540879};
test_output[2143] = '{40.7214903348};
############ END DEBUG ############*/
test_input[17152:17159] = '{32'h4149ad32, 32'h41df909e, 32'h40136ae6, 32'h42aeda72, 32'h428fa592, 32'h42a518f4, 32'hc1dcef79, 32'h42966150};
test_label[2144] = '{32'h42aeda72};
test_output[2144] = '{32'h3bf8ad68};
/*############ DEBUG ############
test_input[17152:17159] = '{12.6047843582, 27.945614217, 2.30339946456, 87.42664744, 71.8233791184, 82.5487341635, -27.6169301654, 75.1900631272};
test_label[2144] = '{87.42664744};
test_output[2144] = '{0.00758903084809};
############ END DEBUG ############*/
test_input[17160:17167] = '{32'hc2938253, 32'h4236111a, 32'h4017132a, 32'h41a3ec10, 32'h424d6fee, 32'hc20eaeca, 32'h42a80835, 32'hc1fe9118};
test_label[2145] = '{32'h4017132a};
test_output[2145] = '{32'h42a34f9c};
/*############ DEBUG ############
test_input[17160:17167] = '{-73.7545400894, 45.5167019769, 2.36054458996, 20.4902641743, 51.3593064679, -35.6706937613, 84.0160288068, -31.8208473643};
test_label[2145] = '{2.36054458996};
test_output[2145] = '{81.6554842168};
############ END DEBUG ############*/
test_input[17168:17175] = '{32'hc14dcd76, 32'h42b2143e, 32'hc29d7e09, 32'h42ab226b, 32'h4234d210, 32'hc1988dab, 32'h41944f17, 32'h424cd252};
test_label[2146] = '{32'hc1988dab};
test_output[2146] = '{32'h42d8474f};
/*############ DEBUG ############
test_input[17168:17175] = '{-12.8626609581, 89.0395318166, -78.7461630826, 85.567223742, 45.2051401358, -19.0691731563, 18.5386181368, 51.2053892051};
test_label[2146] = '{-19.0691731563};
test_output[2146] = '{108.139278108};
############ END DEBUG ############*/
test_input[17176:17183] = '{32'h42501528, 32'h428632d0, 32'h421f5f35, 32'h4107b7c6, 32'hc175da95, 32'h3f333bc3, 32'hc123330e, 32'hc295b3e7};
test_label[2147] = '{32'h3f333bc3};
test_output[2147] = '{32'h4284cc58};
/*############ DEBUG ############
test_input[17176:17183] = '{52.0206620634, 67.0992403335, 39.8429762243, 8.48236636366, -15.3658644666, 0.700130649968, -10.1999643527, -74.8513750371};
test_label[2147] = '{0.700130649968};
test_output[2147] = '{66.3991099663};
############ END DEBUG ############*/
test_input[17184:17191] = '{32'hc26d4bd4, 32'hc1cbd03c, 32'hc1051652, 32'h42262324, 32'h4290d6b0, 32'hc2789990, 32'h429ff755, 32'hc20af9da};
test_label[2148] = '{32'h4290d6b0};
test_output[2148] = '{32'h40f20e84};
/*############ DEBUG ############
test_input[17184:17191] = '{-59.3240506301, -25.4766768019, -8.31794942842, 41.5343157898, 72.4193145058, -62.1499642119, 79.9830674218, -34.7439956337};
test_label[2148] = '{72.4193145058};
test_output[2148] = '{7.56427170554};
############ END DEBUG ############*/
test_input[17192:17199] = '{32'hc2515a4a, 32'hc21fab74, 32'hc2a29d6d, 32'hc2bfc899, 32'h4281a049, 32'hc0a8542a, 32'h4138f2cc, 32'h41f735b0};
test_label[2149] = '{32'h41f735b0};
test_output[2149] = '{32'h4207a5ba};
/*############ DEBUG ############
test_input[17192:17199] = '{-52.3381711793, -39.9174362248, -81.3074730383, -95.8917919261, 64.8130567503, -5.26027379002, 11.5592766601, 30.9012149749};
test_label[2149] = '{30.9012149749};
test_output[2149] = '{33.9118417755};
############ END DEBUG ############*/
test_input[17200:17207] = '{32'h4233fe86, 32'h429e4655, 32'h411ea7db, 32'hc2b000b4, 32'hc2b5f89f, 32'hc21d5bf0, 32'h429c1999, 32'h42766fe3};
test_label[2150] = '{32'h4233fe86};
test_output[2150] = '{32'h4209b79f};
/*############ DEBUG ############
test_input[17200:17207] = '{44.9985578925, 79.1373709204, 9.91598041104, -88.0013706704, -90.9855850159, -39.3397842398, 78.0499958107, 61.6092636528};
test_label[2150] = '{44.9985578925};
test_output[2150] = '{34.4293162737};
############ END DEBUG ############*/
test_input[17208:17215] = '{32'hc07877c4, 32'h4283947b, 32'h424ca3a2, 32'h42c6f42b, 32'hc2ab41fd, 32'hc29820e7, 32'h42bd45c9, 32'hc2a95ff5};
test_label[2151] = '{32'hc2a95ff5};
test_output[2151] = '{32'h43382c14};
/*############ DEBUG ############
test_input[17208:17215] = '{-3.88230997943, 65.78999945, 51.1597967032, 99.4768911866, -85.6288819584, -76.0642658445, 94.6362988233, -84.6874179455};
test_label[2151] = '{-84.6874179455};
test_output[2151] = '{184.172180443};
############ END DEBUG ############*/
test_input[17216:17223] = '{32'h4109a8c8, 32'h425c1c63, 32'h42a3febc, 32'hc14a9382, 32'h421d378d, 32'hc1837f20, 32'h4229548c, 32'hc2aceae7};
test_label[2152] = '{32'hc1837f20};
test_output[2152] = '{32'h42c4de85};
/*############ DEBUG ############
test_input[17216:17223] = '{8.60370603333, 55.0277209706, 81.9975316548, -12.6610129568, 39.3042472488, -16.4370735651, 42.332563776, -86.4587914762};
test_label[2152] = '{-16.4370735651};
test_output[2152] = '{98.4346052199};
############ END DEBUG ############*/
test_input[17224:17231] = '{32'hc10ec033, 32'h403abc9c, 32'h424ce8db, 32'h40ffb600, 32'hc2bb7a5b, 32'h4134ce65, 32'h4288f29f, 32'hc27736e8};
test_label[2153] = '{32'hc2bb7a5b};
test_output[2153] = '{32'h4322367d};
/*############ DEBUG ############
test_input[17224:17231] = '{-8.92192368158, 2.91776170119, 51.227397415, 7.99096670645, -93.7389769173, 11.3003893006, 68.4738690992, -61.8036202666};
test_label[2153] = '{-93.7389769173};
test_output[2153] = '{162.212846049};
############ END DEBUG ############*/
test_input[17232:17239] = '{32'hc2766d5f, 32'hc295270a, 32'hc2ae1ce7, 32'hc282d865, 32'hc2982bb7, 32'h4297c36e, 32'hc11fdad0, 32'hc2531386};
test_label[2154] = '{32'hc2531386};
test_output[2154] = '{32'h4300a699};
/*############ DEBUG ############
test_input[17232:17239] = '{-61.6068061409, -74.5762494076, -87.0564500349, -65.4226430729, -76.0853774902, 75.8816980047, -9.99092116232, -52.7690670218};
test_label[2154] = '{-52.7690670218};
test_output[2154] = '{128.650765026};
############ END DEBUG ############*/
test_input[17240:17247] = '{32'h42c28919, 32'h425c298a, 32'hc048ed4f, 32'hc1871cd6, 32'hc254e271, 32'h417ac833, 32'hc0ccff6a, 32'hc2b0362c};
test_label[2155] = '{32'h417ac833};
test_output[2155] = '{32'h42a33012};
/*############ DEBUG ############
test_input[17240:17247] = '{97.2677670733, 55.0405672278, -3.1394842212, -16.889079188, -53.2211352049, 15.6738763059, -6.40617838898, -88.1058066938};
test_label[2155] = '{15.6738763059};
test_output[2155] = '{81.5938907674};
############ END DEBUG ############*/
test_input[17248:17255] = '{32'hc29e499e, 32'hc194102f, 32'h420d6929, 32'hc27819e7, 32'hc2ad2249, 32'hc29b0481, 32'hc2c2563d, 32'h42c6b7f6};
test_label[2156] = '{32'hc2ad2249};
test_output[2156] = '{32'h4339ed1f};
/*############ DEBUG ############
test_input[17248:17255] = '{-79.1437834724, -18.5079019389, 35.352696165, -62.0252955377, -86.5669603195, -77.508795485, -97.1684315488, 99.3592959467};
test_label[2156] = '{-86.5669603195};
test_output[2156] = '{185.926256266};
############ END DEBUG ############*/
test_input[17256:17263] = '{32'hc22da943, 32'hc2ad3ee9, 32'hc2abbc2c, 32'h426bc085, 32'h428bc0c8, 32'hc2a13a38, 32'h42679ff8, 32'hc17f320f};
test_label[2157] = '{32'hc2a13a38};
test_output[2157] = '{32'h43167d81};
/*############ DEBUG ############
test_input[17256:17263] = '{-43.4152944019, -86.6228734119, -85.8675255702, 58.9380086118, 69.8765258822, -80.6137060659, 57.9062187427, -15.949720992};
test_label[2157] = '{-80.6137060659};
test_output[2157] = '{150.490256038};
############ END DEBUG ############*/
test_input[17264:17271] = '{32'hc2bc5f04, 32'hc24cc1e5, 32'h4227e6d1, 32'hc29a768a, 32'h42340693, 32'h41853276, 32'hc199f84f, 32'hc26c4f16};
test_label[2158] = '{32'hc199f84f};
test_output[2158] = '{32'h42809980};
/*############ DEBUG ############
test_input[17264:17271] = '{-94.1855777782, -51.1893486429, 41.9754049379, -77.2315227461, 45.0064191148, 16.6496382091, -19.2462452312, -59.0772306135};
test_label[2158] = '{-19.2462452312};
test_output[2158] = '{64.2998023483};
############ END DEBUG ############*/
test_input[17272:17279] = '{32'hc195f2cd, 32'hc2c60624, 32'hc128d548, 32'h428f7fad, 32'h42b4cb4f, 32'hc235ff12, 32'hc234aafd, 32'h42901507};
test_label[2159] = '{32'hc2c60624};
test_output[2159] = '{32'h433d68b9};
/*############ DEBUG ############
test_input[17272:17279] = '{-18.7435548165, -99.0119900739, -10.5520701635, 71.7493666037, 90.3970880944, -45.499092299, -45.166980316, 72.0410704971};
test_label[2159] = '{-99.0119900739};
test_output[2159] = '{189.409078187};
############ END DEBUG ############*/
test_input[17280:17287] = '{32'hc1fdc074, 32'h42034b71, 32'hc2769985, 32'hc0bf70bb, 32'hc123c735, 32'h429164ed, 32'hc28f3357, 32'h4261383d};
test_label[2160] = '{32'hc28f3357};
test_output[2160] = '{32'h43104c22};
/*############ DEBUG ############
test_input[17280:17287] = '{-31.7189706136, 32.823673294, -61.6499225971, -5.9825111386, -10.2361342246, 72.6971179787, -71.6002698443, 56.3049189116};
test_label[2160] = '{-71.6002698443};
test_output[2160] = '{144.297387899};
############ END DEBUG ############*/
test_input[17288:17295] = '{32'hc152418d, 32'hc1b49cc5, 32'hc2c1f878, 32'hc23f5f86, 32'h3faa74e3, 32'hc267c538, 32'hc2b11608, 32'h40b2907c};
test_label[2161] = '{32'hc2c1f878};
test_output[2161] = '{32'h42cd28c3};
/*############ DEBUG ############
test_input[17288:17295] = '{-13.1410036954, -22.5765479951, -96.9852903948, -47.8432847209, 1.33169205072, -57.9425975453, -88.543033052, 5.58013721942};
test_label[2161] = '{-96.9852903948};
test_output[2161] = '{102.579612962};
############ END DEBUG ############*/
test_input[17296:17303] = '{32'h4240a87e, 32'hc1b75540, 32'hc2c5fcf9, 32'h42452e64, 32'h403c6793, 32'h42bc8cb3, 32'hc131aca4, 32'h4254fa27};
test_label[2162] = '{32'h403c6793};
test_output[2162] = '{32'h42b6a977};
/*############ DEBUG ############
test_input[17296:17303] = '{48.1645413588, -22.9166264269, -98.9940852936, 49.2953020752, 2.94382168375, 94.2748039363, -11.1046484817, 53.244291267};
test_label[2162] = '{2.94382168375};
test_output[2162] = '{91.3309822526};
############ END DEBUG ############*/
test_input[17304:17311] = '{32'h42624d56, 32'hc27997ba, 32'hc2a83c30, 32'hc2455894, 32'hc2956e47, 32'hc1ab78f6, 32'h429341c4, 32'hc2842925};
test_label[2163] = '{32'hc2a83c30};
test_output[2163] = '{32'h431dbefa};
/*############ DEBUG ############
test_input[17304:17311] = '{56.5755233677, -62.3981719288, -84.1175565126, -49.3365025539, -74.715386338, -21.4340623589, 73.6284506682, -66.0803570038};
test_label[2163] = '{-84.1175565126};
test_output[2163] = '{157.74600722};
############ END DEBUG ############*/
test_input[17312:17319] = '{32'hbee4164d, 32'hc2337075, 32'hc205e483, 32'hc211d573, 32'h41768c31, 32'h418230e5, 32'hc20d6fce, 32'hc1ae72e8};
test_label[2164] = '{32'h418230e5};
test_output[2164] = '{32'h3eb3f80a};
/*############ DEBUG ############
test_input[17312:17319] = '{-0.445482628919, -44.8598195674, -33.4731573196, -36.4584463492, 15.4092264087, 16.2738733965, -35.3591838469, -21.8061068655};
test_label[2164] = '{16.2738733965};
test_output[2164] = '{0.351501775154};
############ END DEBUG ############*/
test_input[17320:17327] = '{32'h41b57b55, 32'h42289ebf, 32'h40daaae6, 32'h4183f412, 32'hc2a6f29e, 32'hc209aea2, 32'hc1b291d3, 32'h4256e23a};
test_label[2165] = '{32'h4183f412};
test_output[2165] = '{32'h4214e833};
/*############ DEBUG ############
test_input[17320:17327] = '{22.6852214034, 42.1550259107, 6.83336184757, 16.49417495, -83.4738602201, -34.4205411713, -22.3212038346, 53.7209228134};
test_label[2165] = '{16.49417495};
test_output[2165] = '{37.2267573475};
############ END DEBUG ############*/
test_input[17328:17335] = '{32'h42b10f96, 32'hc20aa591, 32'hc2bcce10, 32'h41d41930, 32'hc2c3a347, 32'h4245b0f1, 32'h42759b71, 32'h411a8fe0};
test_label[2166] = '{32'hc2bcce10};
test_output[2166] = '{32'h4336eed3};
/*############ DEBUG ############
test_input[17328:17335] = '{88.5304390147, -34.6616843552, -94.4024684077, 26.5122992197, -97.8189031478, 49.4227957391, 61.4017989546, 9.66012562779};
test_label[2166] = '{-94.4024684077};
test_output[2166] = '{182.932907422};
############ END DEBUG ############*/
test_input[17336:17343] = '{32'hc263ed84, 32'h42b90b69, 32'h40e2d128, 32'hc24de12a, 32'h41c9c955, 32'h428740d3, 32'h4249d512, 32'h41ed83d0};
test_label[2167] = '{32'hc24de12a};
test_output[2167] = '{32'h430ffdff};
/*############ DEBUG ############
test_input[17336:17343] = '{-56.981949075, 92.5222860976, 7.08803165281, -51.4698886479, 25.2233060621, 67.6266093452, 50.4580767124, 29.6893624503};
test_label[2167] = '{-51.4698886479};
test_output[2167] = '{143.992174746};
############ END DEBUG ############*/
test_input[17344:17351] = '{32'h4294f62c, 32'hc20cf86f, 32'h40cfae18, 32'hc2880ba4, 32'hc15c7c1b, 32'h4294dc72, 32'h414f280e, 32'hc15fa984};
test_label[2168] = '{32'hc15c7c1b};
test_output[2168] = '{32'h42b1dbe0};
/*############ DEBUG ############
test_input[17344:17351] = '{74.4808065235, -35.2426116152, 6.49000149183, -68.0227378362, -13.7802988458, 74.4305569633, 12.9472790334, -13.9788859022};
test_label[2168] = '{-13.7802988458};
test_output[2168] = '{88.9294433638};
############ END DEBUG ############*/
test_input[17352:17359] = '{32'h405c605d, 32'hbf8f52da, 32'hc2b82a95, 32'hc275c9e9, 32'h42c316ed, 32'hc126601c, 32'hc25cc6f3, 32'h42504a11};
test_label[2169] = '{32'h405c605d};
test_output[2169] = '{32'h42bc33ea};
/*############ DEBUG ############
test_input[17352:17359] = '{3.44338161401, -1.11971591932, -92.0831674244, -61.4471763028, 97.5447744481, -10.39846402, -55.1942867551, 52.0723312142};
test_label[2169] = '{3.44338161401};
test_output[2169] = '{94.1013928341};
############ END DEBUG ############*/
test_input[17360:17367] = '{32'h4280df84, 32'hc28c2edc, 32'h41ca4517, 32'h42129ac9, 32'h40cc47c0, 32'h424c7c9c, 32'hc19f0c87, 32'h42a1e002};
test_label[2170] = '{32'h42129ac9};
test_output[2170] = '{32'h4231253b};
/*############ DEBUG ############
test_input[17360:17367] = '{64.4365535278, -70.0915215366, 25.2837348441, 36.651155978, 6.38375848343, 51.1216898055, -19.8811171174, 80.9375143649};
test_label[2170] = '{36.651155978};
test_output[2170] = '{44.2863584551};
############ END DEBUG ############*/
test_input[17368:17375] = '{32'h40c30ae2, 32'hc29e5b5d, 32'h4259b806, 32'hc2c0ae49, 32'hc29e0bb1, 32'hc212cdb1, 32'h42a91691, 32'hc28551a7};
test_label[2171] = '{32'h4259b806};
test_output[2171] = '{32'h41f0ea3b};
/*############ DEBUG ############
test_input[17368:17375] = '{6.0950783504, -79.1784435309, 54.4297090873, -96.3403987493, -79.0228375685, -36.7008697097, 84.5440786943, -66.6594779};
test_label[2171] = '{54.4297090873};
test_output[2171] = '{30.114369607};
############ END DEBUG ############*/
test_input[17376:17383] = '{32'hc2c16726, 32'hc1f6123d, 32'h42a4d9c8, 32'hc210b17c, 32'h41b088ba, 32'h425c7e55, 32'hc1559db6, 32'hc1da4e14};
test_label[2172] = '{32'hc1559db6};
test_output[2172] = '{32'h42bf8d7f};
/*############ DEBUG ############
test_input[17376:17383] = '{-96.7014609268, -30.7589062865, 82.4253562692, -36.1733237524, 22.0667617643, 55.1233695379, -13.3510038021, -27.2881242965};
test_label[2172] = '{-13.3510038021};
test_output[2172] = '{95.7763600713};
############ END DEBUG ############*/
test_input[17384:17391] = '{32'hc284e56a, 32'h42739fee, 32'h41e73825, 32'h426e91ee, 32'hc1f9fa2b, 32'hc18b1f23, 32'hc25a6619, 32'h429d4231};
test_label[2173] = '{32'h41e73825};
test_output[2173] = '{32'h4246e850};
/*############ DEBUG ############
test_input[17384:17391] = '{-66.4480717301, 60.9061827858, 28.9024142756, 59.6425077991, -31.247152183, -17.3902035123, -54.5997064463, 78.6292830158};
test_label[2173] = '{28.9024142756};
test_output[2173] = '{49.7268687659};
############ END DEBUG ############*/
test_input[17392:17399] = '{32'h428bc7bc, 32'h40eeae39, 32'h4297c2ac, 32'h41bb5aff, 32'h42aa6869, 32'h42993ce8, 32'hc2bfa432, 32'h4256ac96};
test_label[2174] = '{32'h42993ce8};
test_output[2174] = '{32'h41095d29};
/*############ DEBUG ############
test_input[17392:17399] = '{69.89010287, 7.45876763592, 75.8802157466, 23.4194321127, 85.2039276759, 76.6189599034, -95.8206952693, 53.6685411751};
test_label[2174] = '{76.6189599034};
test_output[2174] = '{8.58524413393};
############ END DEBUG ############*/
test_input[17400:17407] = '{32'hc2b3d5b4, 32'h4201129d, 32'hc1839d16, 32'h425b80d2, 32'h421acc5d, 32'hc2b472c7, 32'hc1fe8185, 32'hc11576da};
test_label[2175] = '{32'hc1fe8185};
test_output[2175] = '{32'h42ad60ca};
/*############ DEBUG ############
test_input[17400:17407] = '{-89.9173883827, 32.2681773366, -16.4517012223, 54.8758001834, 38.699573296, -90.224174366, -31.813241264, -9.34151681429};
test_label[2175] = '{-31.813241264};
test_output[2175] = '{86.6890415419};
############ END DEBUG ############*/
test_input[17408:17415] = '{32'hc1ab8764, 32'hc248fea7, 32'h42153155, 32'h42c3dc38, 32'h429fd545, 32'hc2b11afe, 32'h42a4cef4, 32'hc20ba9e3};
test_label[2176] = '{32'h42c3dc38};
test_output[2176] = '{32'h34524210};
/*############ DEBUG ############
test_input[17408:17415] = '{-21.4411082775, -50.2486820687, 37.2981776732, 97.9301134431, 79.9165439571, -88.5527217135, 82.4042024785, -34.9159066771};
test_label[2176] = '{97.9301134431};
test_output[2176] = '{1.95818080605e-07};
############ END DEBUG ############*/
test_input[17416:17423] = '{32'h422349ee, 32'hc27ccc74, 32'h42ba4631, 32'h42a5948f, 32'hc2067117, 32'hc20f9d47, 32'h42be42b9, 32'h428c2da6};
test_label[2177] = '{32'h42be42b9};
test_output[2177] = '{32'h3e02ced6};
/*############ DEBUG ############
test_input[17416:17423] = '{40.8221954734, -63.1996600473, 93.13709609, 82.7901572175, -33.6104401625, -35.9035930107, 95.1303188287, 70.0891565885};
test_label[2177] = '{95.1303188287};
test_output[2177] = '{0.127742144011};
############ END DEBUG ############*/
test_input[17424:17431] = '{32'hc22f502f, 32'hc1b8a6b7, 32'hc0da6160, 32'h42710eb2, 32'h42c2a5b7, 32'h41a1bbab, 32'hc2586e2a, 32'h41331e0d};
test_label[2178] = '{32'h42710eb2};
test_output[2178] = '{32'h42143cbd};
/*############ DEBUG ############
test_input[17424:17431] = '{-43.8283033009, -23.0814043763, -6.82438665983, 60.2643518861, 97.3236652512, 20.2166339873, -54.1075813518, 11.1948362657};
test_label[2178] = '{60.2643518861};
test_output[2178] = '{37.0593133651};
############ END DEBUG ############*/
test_input[17432:17439] = '{32'h41a8aec0, 32'hc2083917, 32'h416f0d4f, 32'hc2a0c347, 32'h41f0dcb7, 32'hc1e6f389, 32'hc2656127, 32'h416d535c};
test_label[2179] = '{32'hc1e6f389};
test_output[2179] = '{32'h426be840};
/*############ DEBUG ############
test_input[17432:17439] = '{21.0853272153, -34.0557506765, 14.9407487987, -80.3814003974, 30.1077708591, -28.8689137004, -57.3448758546, 14.8328517342};
test_label[2179] = '{-28.8689137004};
test_output[2179] = '{58.9768057143};
############ END DEBUG ############*/
test_input[17440:17447] = '{32'hc1c73891, 32'hc1a68edd, 32'hc23bb534, 32'hc2a49d4c, 32'hc2bf96a3, 32'hc1895334, 32'hc2181665, 32'h41071d96};
test_label[2180] = '{32'hc1895334};
test_output[2180] = '{32'h41cce1ff};
/*############ DEBUG ############
test_input[17440:17447] = '{-24.9026200546, -20.8197576009, -46.9269546979, -82.3072208824, -95.7942118024, -17.1656259565, -38.0218702474, 8.44472359708};
test_label[2180] = '{-17.1656259565};
test_output[2180] = '{25.6103495536};
############ END DEBUG ############*/
test_input[17448:17455] = '{32'hc1926037, 32'h422cea85, 32'hc1f9c50f, 32'hc13c61a4, 32'hc2286bf1, 32'hc1a5e15d, 32'hc23630be, 32'h412c02b5};
test_label[2181] = '{32'hc1f9c50f};
test_output[2181] = '{32'h4294e686};
/*############ DEBUG ############
test_input[17448:17455] = '{-18.2969797991, 43.2290217576, -31.221220723, -11.77383792, -42.1054117419, -20.7350403627, -45.5476002588, 10.7506613629};
test_label[2181] = '{-31.221220723};
test_output[2181] = '{74.4502424806};
############ END DEBUG ############*/
test_input[17456:17463] = '{32'hc1994e93, 32'h425e50cd, 32'hc1eeff98, 32'hc29f38df, 32'hc2988b04, 32'h420cb167, 32'h412533f7, 32'h426e2377};
test_label[2182] = '{32'hc1994e93};
test_output[2182] = '{32'h429d6f16};
/*############ DEBUG ############
test_input[17456:17463] = '{-19.1633663916, 55.5789078438, -29.874801268, -79.6110767961, -76.2715152935, 35.1732441603, 10.3251868514, 59.5346351394};
test_label[2182] = '{-19.1633663916};
test_output[2182] = '{78.716965316};
############ END DEBUG ############*/
test_input[17464:17471] = '{32'h421450f4, 32'hc11777aa, 32'h408e5287, 32'hc29b1cc4, 32'hc2728c6d, 32'h428d081d, 32'hc1ff318a, 32'hc29e58aa};
test_label[2183] = '{32'h408e5287};
test_output[2183] = '{32'h428422f4};
/*############ DEBUG ############
test_input[17464:17471] = '{37.0790550926, -9.46671473183, 4.4475741898, -77.5561846868, -60.6371363622, 70.5158444158, -31.8991885269, -79.1731710716};
test_label[2183] = '{4.4475741898};
test_output[2183] = '{66.068270226};
############ END DEBUG ############*/
test_input[17472:17479] = '{32'h422992b4, 32'h42bd200a, 32'h42a5a946, 32'hc2aee88d, 32'hc2bad415, 32'h429a795f, 32'h42977c9e, 32'hc1b4ed91};
test_label[2184] = '{32'h42977c9e};
test_output[2184] = '{32'h41968db6};
/*############ DEBUG ############
test_input[17472:17479] = '{42.3932646445, 94.5625798527, 82.8306149356, -87.4542035642, -93.4142206202, 77.2370561797, 75.7433922055, -22.6159986024};
test_label[2184] = '{75.7433922055};
test_output[2184] = '{18.8191957166};
############ END DEBUG ############*/
test_input[17480:17487] = '{32'hc2c5c788, 32'h42a32cc1, 32'hc230321f, 32'h42b44d4e, 32'hc1a558c7, 32'h4142495f, 32'h429b0641, 32'hc1568503};
test_label[2185] = '{32'hc2c5c788};
test_output[2185] = '{32'h433d0a77};
/*############ DEBUG ############
test_input[17480:17487] = '{-98.8897061413, 81.5874092577, -44.0489476826, 90.1509840669, -20.6683492513, 12.142912812, 77.5122165447, -13.4074731498};
test_label[2185] = '{-98.8897061413};
test_output[2185] = '{189.040884369};
############ END DEBUG ############*/
test_input[17488:17495] = '{32'h42438188, 32'h41570077, 32'h4230fee5, 32'h42c31c89, 32'hc1cc61fc, 32'h416bb8f8, 32'h41edb319, 32'h41ecdc62};
test_label[2186] = '{32'h416bb8f8};
test_output[2186] = '{32'h42a5a56a};
/*############ DEBUG ############
test_input[17488:17495] = '{48.8764964282, 13.4376134595, 44.2489198888, 97.555733857, -25.547843377, 14.7326586458, 29.7124497203, 29.6076097299};
test_label[2186] = '{14.7326586458};
test_output[2186] = '{82.8230752112};
############ END DEBUG ############*/
test_input[17496:17503] = '{32'h4296ed2f, 32'h411d0bc0, 32'hc2acef3a, 32'hc2b0ba85, 32'hc1016f0a, 32'hc1a9225a, 32'h423d2cda, 32'h3ec6ed38};
test_label[2187] = '{32'hc2acef3a};
test_output[2187] = '{32'h4321ee34};
/*############ DEBUG ############
test_input[17496:17503] = '{75.4632473939, 9.81536860837, -86.4672410746, -88.364293232, -8.08960952827, -21.1417727051, 47.2937990315, 0.388528591581};
test_label[2187] = '{-86.4672410746};
test_output[2187] = '{161.930488469};
############ END DEBUG ############*/
test_input[17504:17511] = '{32'hc217f035, 32'hc13fa6a3, 32'h42c3ce19, 32'h428702c7, 32'hc25e8183, 32'hc2a1afd8, 32'h429d63c2, 32'h411ff9de};
test_label[2188] = '{32'hc217f035};
test_output[2188] = '{32'h4307e31a};
/*############ DEBUG ############
test_input[17504:17511] = '{-37.9845767175, -11.9781825285, 97.9025311478, 67.5054226859, -55.6264751107, -80.8434455363, 78.6948394919, 9.99850258327};
test_label[2188] = '{-37.9845767175};
test_output[2188] = '{135.88710787};
############ END DEBUG ############*/
test_input[17512:17519] = '{32'h424049e7, 32'hc283d02d, 32'hc0dcce29, 32'h42977c75, 32'h4257672e, 32'hc295bfbf, 32'h42bc2c21, 32'h41b60227};
test_label[2189] = '{32'h42977c75};
test_output[2189] = '{32'h4192beae};
/*############ DEBUG ############
test_input[17512:17519] = '{48.0721710219, -65.9065923435, -6.9001659004, 75.7430825138, 53.8507617494, -74.8745028706, 94.0861884452, 22.7510518035};
test_label[2189] = '{75.7430825138};
test_output[2189] = '{18.3431059422};
############ END DEBUG ############*/
test_input[17520:17527] = '{32'h4222f4a7, 32'h42458b0b, 32'hc0fd7a2d, 32'hc1da56f1, 32'h4232fc75, 32'h4210e092, 32'h41f1ec45, 32'h41f5691b};
test_label[2190] = '{32'h4232fc75};
test_output[2190] = '{32'h4094c4ef};
/*############ DEBUG ############
test_input[17520:17527] = '{40.7389192407, 49.3857854853, -7.92116400937, -27.2924524055, 44.7465402275, 36.2193069049, 30.2403664244, 30.6763209846};
test_label[2190] = '{44.7465402275};
test_output[2190] = '{4.649039727};
############ END DEBUG ############*/
test_input[17528:17535] = '{32'h42b4be61, 32'hc294d38e, 32'hc2acaaf3, 32'h40ec93da, 32'h42428aad, 32'h422e9eb8, 32'hc2041ece, 32'h4192b0b3};
test_label[2191] = '{32'h42428aad};
test_output[2191] = '{32'h4226f215};
/*############ DEBUG ############
test_input[17528:17535] = '{90.3718362443, -74.4131933351, -86.3338835692, 7.39304826675, 48.6354263554, 43.6549976956, -33.0300820893, 18.3362791482};
test_label[2191] = '{48.6354263554};
test_output[2191] = '{41.7364098889};
############ END DEBUG ############*/
test_input[17536:17543] = '{32'hc29b573f, 32'h414beecc, 32'hc28128ba, 32'hc057d850, 32'hc2964185, 32'h42578af7, 32'hc197c5d1, 32'h410d92b0};
test_label[2192] = '{32'hc29b573f};
test_output[2192] = '{32'h43038e5d};
/*############ DEBUG ############
test_input[17536:17543] = '{-77.6704007675, 12.7457997571, -64.5795458344, -3.37257756583, -75.1279683787, 53.8857081563, -18.9715895267, 8.84831275593};
test_label[2192] = '{-77.6704007675};
test_output[2192] = '{131.556108924};
############ END DEBUG ############*/
test_input[17544:17551] = '{32'hc2b8bd74, 32'hc28388fd, 32'hc22d5f5e, 32'hc0fea35e, 32'h428808fa, 32'h421f1af8, 32'hc1b45462, 32'h42b0d3de};
test_label[2193] = '{32'hc28388fd};
test_output[2193] = '{32'h431a2e6e};
/*############ DEBUG ############
test_input[17544:17551] = '{-92.3700281177, -65.7675557021, -43.3431336666, -7.95744228728, 68.0175333953, 39.7763353933, -22.5412020239, 88.41380467};
test_label[2193] = '{-65.7675557021};
test_output[2193] = '{154.181360374};
############ END DEBUG ############*/
test_input[17552:17559] = '{32'h4223629f, 32'h42466f7e, 32'hc27643ae, 32'hc2a8d1db, 32'h427fcb0f, 32'h41240df6, 32'hbfedce5f, 32'hc29e644c};
test_label[2194] = '{32'h4223629f};
test_output[2194] = '{32'h41b8d0df};
/*############ DEBUG ############
test_input[17552:17559] = '{40.846310783, 49.6088798862, -61.5660928695, -84.4098709893, 63.9482981166, 10.2534084231, -1.85786045827, -79.195888681};
test_label[2194] = '{40.846310783};
test_output[2194] = '{23.1019879259};
############ END DEBUG ############*/
test_input[17560:17567] = '{32'h422ce698, 32'hc21a1ec4, 32'h42c1f76e, 32'hc1d79885, 32'h4001fa17, 32'hc29f4c76, 32'hc27e5539, 32'hbfce5f3b};
test_label[2195] = '{32'hc21a1ec4};
test_output[2195] = '{32'h43078368};
/*############ DEBUG ############
test_input[17560:17567] = '{43.2251876252, -38.5300431784, 96.9832582993, -26.9494723045, 2.03088936544, -79.6493361091, -63.5832235379, -1.61228116212};
test_label[2195] = '{-38.5300431784};
test_output[2195] = '{135.513301478};
############ END DEBUG ############*/
test_input[17568:17575] = '{32'hc2b8e8aa, 32'hc2b8e643, 32'hc2a8f7bb, 32'h42a2d798, 32'hc21ac608, 32'h4263096f, 32'hc2a9557f, 32'h42c6fab4};
test_label[2196] = '{32'h42c6fab4};
test_output[2196] = '{32'h32744f14};
/*############ DEBUG ############
test_input[17568:17575] = '{-92.454423859, -92.4497276451, -84.4838490779, 81.4210846363, -38.6933884183, 56.7592112963, -84.6669868641, 99.4896553372};
test_label[2196] = '{99.4896553372};
test_output[2196] = '{1.422064987e-08};
############ END DEBUG ############*/
test_input[17576:17583] = '{32'hc2a6c376, 32'h42bf9395, 32'h4282e4f3, 32'hc27bdb0c, 32'h4189bb63, 32'h42267071, 32'hc2b80070, 32'hc2bee99f};
test_label[2197] = '{32'hc2bee99f};
test_output[2197] = '{32'h433f3e9a};
/*############ DEBUG ############
test_input[17576:17583] = '{-83.3817594992, 95.7882429364, 65.4471686343, -62.9639140857, 17.2164977072, 41.6098050513, -92.0008531305, -95.4562941331};
test_label[2197] = '{-95.4562941331};
test_output[2197] = '{191.24453707};
############ END DEBUG ############*/
test_input[17584:17591] = '{32'h428f0a5f, 32'hc2b8cfa7, 32'h41b06e43, 32'h42555f22, 32'h42c786eb, 32'hc1bdf268, 32'h4294af06, 32'h427e6e44};
test_label[2198] = '{32'h4294af06};
test_output[2198] = '{32'h41cb5f92};
/*############ DEBUG ############
test_input[17584:17591] = '{71.52025855, -92.4055745446, 22.0538378294, 53.3429049296, 99.7635098466, -23.7433624081, 74.3418437929, 63.607679713};
test_label[2198] = '{74.3418437929};
test_output[2198] = '{25.4216660537};
############ END DEBUG ############*/
test_input[17592:17599] = '{32'hc0bdffc1, 32'h401ef2b3, 32'h42b6a0d3, 32'h42c4382d, 32'hc008ddfb, 32'h4288a62b, 32'hc21a664a, 32'h41a84d73};
test_label[2199] = '{32'h42b6a0d3};
test_output[2199] = '{32'h40d97ec1};
/*############ DEBUG ############
test_input[17592:17599] = '{-5.93746992479, 2.48356311559, 91.314111706, 98.1097164769, -2.1385486931, 68.3245495983, -38.5998926253, 21.0378168539};
test_label[2199] = '{91.314111706};
test_output[2199] = '{6.7967228269};
############ END DEBUG ############*/
test_input[17600:17607] = '{32'h4133aff5, 32'hc2612de6, 32'hc2ad2ce7, 32'h427252d3, 32'hc2c2e7fa, 32'hc21620ef, 32'hc292727f, 32'h403431c6};
test_label[2200] = '{32'hc292727f};
test_output[2200] = '{32'h4305cdf4};
/*############ DEBUG ############
test_input[17600:17607] = '{11.2304578934, -56.2948232308, -86.5876963984, 60.5808837066, -97.4530763323, -37.5321632164, -73.2236230224, 2.81553782834};
test_label[2200] = '{-73.2236230224};
test_output[2200] = '{133.804506729};
############ END DEBUG ############*/
test_input[17608:17615] = '{32'hc2a1a388, 32'hc259bb06, 32'h4242b159, 32'hc1a1b83b, 32'hbff079ab, 32'hc2bb7f87, 32'hc1a3f0bd, 32'hc2a89bfb};
test_label[2201] = '{32'hc1a1b83b};
test_output[2201] = '{32'h4289c6bb};
/*############ DEBUG ############
test_input[17608:17615] = '{-80.8193972345, -54.4326397194, 48.6731894675, -20.2149556119, -1.8787129757, -93.7490754178, -20.4925480746, -84.3046479251};
test_label[2201] = '{-20.2149556119};
test_output[2201] = '{68.8881450793};
############ END DEBUG ############*/
test_input[17616:17623] = '{32'h4292948a, 32'h41f91bba, 32'h420a48e6, 32'h41b8fd21, 32'h41843400, 32'hc2c30d39, 32'h42235743, 32'hc297c394};
test_label[2202] = '{32'h41843400};
test_output[2202] = '{32'h42630f15};
/*############ DEBUG ############
test_input[17616:17623] = '{73.2901181019, 31.1385378427, 34.5711898667, 23.1235988039, 16.5253901127, -97.5258220112, 40.8352178602, -75.8819906362};
test_label[2202] = '{16.5253901127};
test_output[2202] = '{56.7647279892};
############ END DEBUG ############*/
test_input[17624:17631] = '{32'hc2abd841, 32'hc2c07bb2, 32'hc2ac8bd7, 32'hc28b0fa4, 32'hc1f81627, 32'h41d81ccc, 32'h42550f41, 32'h3fdf49c4};
test_label[2203] = '{32'hc28b0fa4};
test_output[2203] = '{32'h42f59745};
/*############ DEBUG ############
test_input[17624:17631] = '{-85.9223738364, -96.2415940623, -86.2731230449, -69.5305477359, -31.0108167531, 27.0140603856, 53.2648971566, 1.74443862638};
test_label[2203] = '{-69.5305477359};
test_output[2203] = '{122.795444893};
############ END DEBUG ############*/
test_input[17632:17639] = '{32'hc27166f9, 32'h42036a44, 32'h42892822, 32'hc2a3b855, 32'hc121f9b8, 32'hc2c6c952, 32'h42a04b63, 32'h42a9ffe1};
test_label[2204] = '{32'hc2c6c952};
test_output[2204] = '{32'h43386697};
/*############ DEBUG ############
test_input[17632:17639] = '{-60.3505575765, 32.8537742339, 68.5783822908, -81.8600204297, -10.1234667364, -99.3932072319, 80.1472388489, 84.999761833};
test_label[2204] = '{-99.3932072319};
test_output[2204] = '{184.40074746};
############ END DEBUG ############*/
test_input[17640:17647] = '{32'hc2bce2c4, 32'h425bcde6, 32'h424ef522, 32'h42a58ad7, 32'h42bab2e8, 32'h4241d87b, 32'hc2bd41a8, 32'h418c7722};
test_label[2205] = '{32'h4241d87b};
test_output[2205] = '{32'h42338d5b};
/*############ DEBUG ############
test_input[17640:17647] = '{-94.4429049166, 54.9510743303, 51.7393887975, 82.7711690867, 93.3494233675, 48.4614067223, -94.6282373482, 17.5581704395};
test_label[2205] = '{48.4614067223};
test_output[2205] = '{44.8880421087};
############ END DEBUG ############*/
test_input[17648:17655] = '{32'hc1663a32, 32'hc2af8509, 32'hc246142e, 32'h42a13722, 32'hc29447d4, 32'hc2c38805, 32'hc262016a, 32'hc2c682e5};
test_label[2206] = '{32'hc2af8509};
test_output[2206] = '{32'h43285e16};
/*############ DEBUG ############
test_input[17648:17655] = '{-14.3892078444, -87.7598335017, -49.5197048791, 80.6076845776, -74.1402877556, -97.7656636629, -56.5013826831, -99.2556512546};
test_label[2206] = '{-87.7598335017};
test_output[2206] = '{168.367518079};
############ END DEBUG ############*/
test_input[17656:17663] = '{32'h424214fd, 32'hc226b036, 32'hc1db0c31, 32'h3ff9a93d, 32'hc1b79b35, 32'hc0d99870, 32'h4255f420, 32'h426ec272};
test_label[2207] = '{32'h426ec272};
test_output[2207] = '{32'h3b059759};
/*############ DEBUG ############
test_input[17656:17663] = '{48.5204960273, -41.6720792372, -27.3809533759, 1.95047725562, -22.9507851867, -6.79985823183, 53.4884018335, 59.6898865553};
test_label[2207] = '{59.6898865553};
test_output[2207] = '{0.00203843992884};
############ END DEBUG ############*/
test_input[17664:17671] = '{32'hc2b3e4e9, 32'hc288c39e, 32'h422334b8, 32'h4294149d, 32'h4255c913, 32'h4196224d, 32'h42a94253, 32'h422c2a8d};
test_label[2208] = '{32'h4255c913};
test_output[2208] = '{32'h41f97735};
/*############ DEBUG ############
test_input[17664:17671] = '{-89.9470889362, -68.3820672881, 40.8014823737, 74.0402640952, 53.4463620961, 18.766749168, 84.6295430896, 43.0415545188};
test_label[2208] = '{53.4463620961};
test_output[2208] = '{31.1832061778};
############ END DEBUG ############*/
test_input[17672:17679] = '{32'hc2bdc320, 32'h42b891bc, 32'hc2703749, 32'hc2c1f49a, 32'hc2356d83, 32'h42351164, 32'h41c10135, 32'h4268a13d};
test_label[2209] = '{32'h41c10135};
test_output[2209] = '{32'h4288516e};
/*############ DEBUG ############
test_input[17672:17679] = '{-94.8811054004, 92.2846354631, -60.0539896645, -96.9777362859, -45.356945232, 45.2669833947, 24.1255898539, 58.1574600869};
test_label[2209] = '{24.1255898539};
test_output[2209] = '{68.1590456092};
############ END DEBUG ############*/
test_input[17680:17687] = '{32'hc2bbb4f7, 32'h424006bc, 32'h42bf0d57, 32'hc1f7a706, 32'hc1f99cb1, 32'h42a13b22, 32'hc0b55359, 32'hc2c42cc9};
test_label[2210] = '{32'hc2c42cc9};
test_output[2210] = '{32'h43419d10};
/*############ DEBUG ############
test_input[17680:17687] = '{-93.8534467121, 48.0065773018, 95.5260545937, -30.9565534829, -31.2015090768, 80.6154925096, -5.66642416308, -98.0874741098};
test_label[2210] = '{-98.0874741098};
test_output[2210] = '{193.613529038};
############ END DEBUG ############*/
test_input[17688:17695] = '{32'hc2ba799e, 32'h41a03ad2, 32'hc2704d6a, 32'h427dba80, 32'h42195d3f, 32'h4163c25f, 32'hc23853a7, 32'hc1bb1630};
test_label[2211] = '{32'h41a03ad2};
test_output[2211] = '{32'h422d9d17};
/*############ DEBUG ############
test_input[17688:17695] = '{-93.2375304487, 20.0287205679, -60.0756002863, 63.4321278043, 38.3410624075, 14.2349541655, -46.0816918788, -23.38583316};
test_label[2211] = '{20.0287205679};
test_output[2211] = '{43.4034072364};
############ END DEBUG ############*/
test_input[17696:17703] = '{32'hc28b5774, 32'h412ddfa4, 32'h423711a9, 32'hc1e51b0c, 32'h428f4466, 32'h42ac6173, 32'hc2981266, 32'hc29302fe};
test_label[2212] = '{32'h428f4466};
test_output[2212] = '{32'h4168e86c};
/*############ DEBUG ############
test_input[17696:17703] = '{-69.6708069327, 10.8670994109, 45.767245218, -28.6382061871, 71.6335872188, 86.1903302653, -76.0359376129, -73.5058471054};
test_label[2212] = '{71.6335872188};
test_output[2212] = '{14.5567435231};
############ END DEBUG ############*/
test_input[17704:17711] = '{32'hc2462dce, 32'h428e17f4, 32'h4241e73c, 32'h42154bc9, 32'h42ab47a0, 32'hc15d1aad, 32'hc2991a31, 32'hc23e36ee};
test_label[2213] = '{32'hc2991a31};
test_output[2213] = '{32'h432230e9};
/*############ DEBUG ############
test_input[17704:17711] = '{-49.5447292691, 71.0467830611, 48.4758142109, 37.3240097848, 85.6398960883, -13.8190130927, -76.5511524571, -47.5536438825};
test_label[2213] = '{-76.5511524571};
test_output[2213] = '{162.191049005};
############ END DEBUG ############*/
test_input[17712:17719] = '{32'hc2b5cc8c, 32'hc2b9d587, 32'hc2c2d305, 32'hc215e936, 32'h42a9a5f6, 32'h42aced93, 32'h4214d24e, 32'h42bffcf5};
test_label[2214] = '{32'hc2c2d305};
test_output[2214] = '{32'h43416803};
/*############ DEBUG ############
test_input[17712:17719] = '{-90.8995068054, -92.9170482277, -97.4121460108, -37.4777466, 84.8241414231, 86.464012725, 37.2053761002, 95.9940559284};
test_label[2214] = '{-97.4121460108};
test_output[2214] = '{193.406288664};
############ END DEBUG ############*/
test_input[17720:17727] = '{32'h429c6f0b, 32'h42c512ee, 32'hc1f13b99, 32'hc222d445, 32'hc2c3c510, 32'hc24e4383, 32'hc2428cbf, 32'hc2be6192};
test_label[2215] = '{32'hc24e4383};
test_output[2215] = '{32'h43161a58};
/*############ DEBUG ############
test_input[17720:17727] = '{78.2168805675, 98.5369710146, -30.1540997499, -40.7072962837, -97.8848844508, -51.5659304925, -48.6374481939, -95.1905675137};
test_label[2215] = '{-51.5659304925};
test_output[2215] = '{150.102901509};
############ END DEBUG ############*/
test_input[17728:17735] = '{32'h42a70277, 32'hc2818df7, 32'hc29b3118, 32'hc16ef0bb, 32'h41f99b26, 32'h4209867d, 32'hc2811c59, 32'h41cf2b34};
test_label[2216] = '{32'h42a70277};
test_output[2216] = '{32'h80000000};
/*############ DEBUG ############
test_input[17728:17735] = '{83.5048117663, -64.7772730766, -77.5958865776, -14.9337718208, 31.2007558157, 34.3813376552, -64.5553632363, 25.8960945016};
test_label[2216] = '{83.5048117663};
test_output[2216] = '{-0.0};
############ END DEBUG ############*/
test_input[17736:17743] = '{32'hc142467e, 32'hc2166e62, 32'hc2c0ec9b, 32'h42144e6a, 32'h421e4d5a, 32'h42268c33, 32'h420b93ed, 32'hc2aad68e};
test_label[2217] = '{32'h42268c33};
test_output[2217] = '{32'h3e05331a};
/*############ DEBUG ############
test_input[17736:17743] = '{-12.1422100968, -37.6077942258, -96.4621187406, 37.076577182, 39.5755380993, 41.636914603, 34.8944596168, -85.4190514348};
test_label[2217] = '{41.636914603};
test_output[2217] = '{0.13007774631};
############ END DEBUG ############*/
test_input[17744:17751] = '{32'h416c952d, 32'h4192e521, 32'hc21dff5f, 32'hc29bf233, 32'h424285fc, 32'hc23ce528, 32'h42abd7ee, 32'hc21f68e5};
test_label[2218] = '{32'hc23ce528};
test_output[2218] = '{32'h43052541};
/*############ DEBUG ############
test_input[17744:17751] = '{14.7864201352, 18.36187911, -39.4993865791, -77.9730417307, 48.6308448386, -47.2237870482, 85.9217406171, -39.8524360042};
test_label[2218] = '{-47.2237870482};
test_output[2218] = '{133.145527665};
############ END DEBUG ############*/
test_input[17752:17759] = '{32'hc2bc3123, 32'hc2ae90f3, 32'h42330f4f, 32'h42b48cb7, 32'h4218f704, 32'hc1fa9c69, 32'hc2855d85, 32'hc2b32c53};
test_label[2219] = '{32'h4218f704};
test_output[2219] = '{32'h4250226a};
/*############ DEBUG ############
test_input[17752:17759] = '{-94.0959698009, -87.2831015781, 44.7649479768, 90.2748347201, 38.2412263068, -31.3263713976, -66.6826565423, -89.5865707463};
test_label[2219] = '{38.2412263068};
test_output[2219] = '{52.0336084133};
############ END DEBUG ############*/
test_input[17760:17767] = '{32'hc06f6ce8, 32'hc1e11392, 32'h42a7d6d7, 32'hc24d84b6, 32'hc2b04afe, 32'hc283768e, 32'h4060b4f9, 32'h42bdf057};
test_label[2220] = '{32'h4060b4f9};
test_output[2220] = '{32'h42b6eab1};
/*############ DEBUG ############
test_input[17760:17767] = '{-3.74102207964, -28.134555162, 83.9196092027, -51.3796020064, -88.1464655264, -65.7315545316, 3.51104578866, 94.969414115};
test_label[2220] = '{3.51104578866};
test_output[2220] = '{91.4583842165};
############ END DEBUG ############*/
test_input[17768:17775] = '{32'h41aef211, 32'h41ad6e3a, 32'h42b52e8e, 32'h4206c3a5, 32'h41d0dc06, 32'h42923cbc, 32'hc29f6e8e, 32'h4171b5b2};
test_label[2221] = '{32'h41d0dc06};
test_output[2221] = '{32'h4280f78c};
/*############ DEBUG ############
test_input[17768:17775] = '{21.8681961836, 21.6788209534, 90.5909264727, 33.6910584846, 26.1074341598, 73.1186186816, -79.715928868, 15.1068589054};
test_label[2221] = '{26.1074341598};
test_output[2221] = '{64.4834923388};
############ END DEBUG ############*/
test_input[17776:17783] = '{32'h4104e350, 32'hc1c60a52, 32'h42b94e93, 32'hc207007a, 32'h4290a4f2, 32'h41607d8a, 32'h412c82d1, 32'h423a0c69};
test_label[2222] = '{32'h412c82d1};
test_output[2222] = '{32'h42a3be39};
/*############ DEBUG ############
test_input[17776:17783] = '{8.30549620461, -24.7550400452, 92.6534685123, -33.7504642562, 72.3221586093, 14.0306491298, 10.7819375426, 46.5121197632};
test_label[2222] = '{10.7819375426};
test_output[2222] = '{81.8715309711};
############ END DEBUG ############*/
test_input[17784:17791] = '{32'hc2aa1ff0, 32'h428aa672, 32'hc2a82828, 32'h423b1a2e, 32'h42c3aeb1, 32'h4243b59d, 32'hc1ac64c3, 32'hc1b6ecda};
test_label[2223] = '{32'h4243b59d};
test_output[2223] = '{32'h4243a7c5};
/*############ DEBUG ############
test_input[17784:17791] = '{-85.0623780722, 69.3250884191, -84.0784294091, 46.7755662334, 97.8411915506, 48.9273549997, -21.5492009992, -22.8656504268};
test_label[2223] = '{48.9273549997};
test_output[2223] = '{48.9138365509};
############ END DEBUG ############*/
test_input[17792:17799] = '{32'hc2b436b4, 32'h4222c396, 32'h42c5b1e0, 32'hc290b924, 32'hc2a38baa, 32'h42a45171, 32'h4283943c, 32'hc21eb0b3};
test_label[2224] = '{32'hc2a38baa};
test_output[2224] = '{32'h43349ec5};
/*############ DEBUG ############
test_input[17792:17799] = '{-90.1068412152, 40.6910026361, 98.847413302, -72.3616026165, -81.7727840634, 82.1590625034, 65.7895239449, -39.6725582195};
test_label[2224] = '{-81.7727840634};
test_output[2224] = '{180.620197422};
############ END DEBUG ############*/
test_input[17800:17807] = '{32'hc179227c, 32'hc15d6389, 32'h42b3ddee, 32'h42c15ed3, 32'hc2bdb0f2, 32'hc1d66aac, 32'hc2a6a53b, 32'hc261597c};
test_label[2225] = '{32'hc1d66aac};
test_output[2225] = '{32'h42f6fa17};
/*############ DEBUG ############
test_input[17800:17807] = '{-15.5709185865, -13.8368007462, 89.9334561144, 96.6852045135, -94.8455982046, -26.8020861569, -83.3227182041, -56.3373852731};
test_label[2225] = '{-26.8020861569};
test_output[2225] = '{123.488458822};
############ END DEBUG ############*/
test_input[17808:17815] = '{32'h4243015d, 32'h42a74ab1, 32'h421b3be7, 32'h4290424c, 32'h428b31d6, 32'hc10ee2fe, 32'hc2b3a715, 32'h4293433a};
test_label[2226] = '{32'h42a74ab1};
test_output[2226] = '{32'h3868c6f5};
/*############ DEBUG ############
test_input[17808:17815] = '{48.7513314995, 83.6458853344, 38.80849875, 72.1294823228, 69.5973381739, -8.93041812743, -89.8263296639, 73.6312993983};
test_label[2226] = '{83.6458853344};
test_output[2226] = '{5.54984047467e-05};
############ END DEBUG ############*/
test_input[17816:17823] = '{32'hc0bb2159, 32'h42bd041e, 32'h4282d33c, 32'hc167dca2, 32'hc271e2ee, 32'h42833746, 32'h40b37126, 32'h40eb94f5};
test_label[2227] = '{32'h40b37126};
test_output[2227] = '{32'h42b1cd0b};
/*############ DEBUG ############
test_input[17816:17823] = '{-5.84782062847, 94.508038217, 65.4125654758, -14.4913650914, -60.4716124568, 65.6079561943, 5.60756207853, 7.36193321633};
test_label[2227] = '{5.60756207853};
test_output[2227] = '{88.9004761385};
############ END DEBUG ############*/
test_input[17824:17831] = '{32'hc1f7f78e, 32'h421d1858, 32'h40d2ff43, 32'hc18f8a35, 32'hc29b0318, 32'h422fed0a, 32'hc2978f13, 32'h4292813a};
test_label[2228] = '{32'h422fed0a};
test_output[2228] = '{32'h41ea2ad3};
/*############ DEBUG ############
test_input[17824:17831] = '{-30.9958772057, 39.2737726997, 6.59366008846, -17.94248426, -77.5060448202, 43.9814816142, -75.7794386585, 73.2523925005};
test_label[2228] = '{43.9814816142};
test_output[2228] = '{29.2709108863};
############ END DEBUG ############*/
test_input[17832:17839] = '{32'hc27f685a, 32'h41071bb2, 32'hc18cf070, 32'hc0dc4379, 32'h424d89a9, 32'h42888ef7, 32'hc299b7e0, 32'h422d9853};
test_label[2229] = '{32'h424d89a9};
test_output[2229] = '{32'h4187288c};
/*############ DEBUG ############
test_input[17832:17839] = '{-63.8519071744, 8.44426198732, -17.6174013201, -6.88323629256, 51.3844345149, 68.279231888, -76.859134288, 43.3987542333};
test_label[2229] = '{51.3844345149};
test_output[2229] = '{16.8947974192};
############ END DEBUG ############*/
test_input[17840:17847] = '{32'hc273f99d, 32'hc20a3b59, 32'h4240cbac, 32'h4226a371, 32'h42c37b11, 32'h41b5122b, 32'hc28b051c, 32'h4233ae44};
test_label[2230] = '{32'h4240cbac};
test_output[2230] = '{32'h42462a77};
/*############ DEBUG ############
test_input[17840:17847] = '{-60.9937614493, -34.5579583464, 48.1988985518, 41.6596122943, 97.7403668803, 22.633870802, -69.5099761615, 44.9201820779};
test_label[2230] = '{48.1988985518};
test_output[2230] = '{49.5414683285};
############ END DEBUG ############*/
test_input[17848:17855] = '{32'h4239f63a, 32'h4266601f, 32'h40213765, 32'hc1f285bb, 32'h428a3b55, 32'h42a10549, 32'hc23e2091, 32'h405332a1};
test_label[2231] = '{32'h405332a1};
test_output[2231] = '{32'h429a6bb5};
/*############ DEBUG ############
test_input[17848:17855] = '{46.4904557097, 57.5938674955, 2.51900606066, -30.3152982108, 69.115881113, 80.5103207682, -47.5318048674, 3.29996516562};
test_label[2231] = '{3.29996516562};
test_output[2231] = '{77.2103668606};
############ END DEBUG ############*/
test_input[17856:17863] = '{32'h42310a13, 32'hc289e0df, 32'h4290b4e0, 32'h426da470, 32'hc2970ee9, 32'hc11a7ea5, 32'hc21ec0b9, 32'h4288ff14};
test_label[2232] = '{32'hc11a7ea5};
test_output[2232] = '{32'h42a40f6f};
/*############ DEBUG ############
test_input[17856:17863] = '{44.2598397767, -68.9392045663, 72.3532677818, 59.4105845406, -75.5291200653, -9.65591906586, -39.6882066442, 68.4981967909};
test_label[2232] = '{-9.65591906586};
test_output[2232] = '{82.0301402771};
############ END DEBUG ############*/
test_input[17864:17871] = '{32'h426a5627, 32'h424df55e, 32'hc1c7e17f, 32'hc2775689, 32'h41422a32, 32'hc28d2d64, 32'hc27325b8, 32'h429009c8};
test_label[2233] = '{32'hc28d2d64};
test_output[2233] = '{32'h430e9b96};
/*############ DEBUG ############
test_input[17864:17871] = '{58.584133116, 51.4896146736, -24.9851055146, -61.8345063813, 12.1353013236, -70.5886563485, -60.7868339937, 72.0191008984};
test_label[2233] = '{-70.5886563485};
test_output[2233] = '{142.607758711};
############ END DEBUG ############*/
test_input[17872:17879] = '{32'h42134f68, 32'hc20f8551, 32'h425869d1, 32'h41983739, 32'hc26b97f2, 32'h42c207c6, 32'h42434715, 32'h429c8ced};
test_label[2234] = '{32'h41983739};
test_output[2234] = '{32'h429bf9f8};
/*############ DEBUG ############
test_input[17872:17879] = '{36.8275440681, -35.8801903425, 54.103335795, 19.0269640383, -58.8983847441, 97.0151829709, 48.8194167284, 78.2752470644};
test_label[2234] = '{19.0269640383};
test_output[2234] = '{77.9882189399};
############ END DEBUG ############*/
test_input[17880:17887] = '{32'hc256cdcc, 32'h403b9e50, 32'h42bbc9e2, 32'hc2572a88, 32'h429bb004, 32'h41d6a3cd, 32'h420c0009, 32'h420fdc44};
test_label[2235] = '{32'h420fdc44};
test_output[2235] = '{32'h4267b780};
/*############ DEBUG ############
test_input[17880:17887] = '{-53.700972222, 2.93153757447, 93.8943027607, -53.7915358523, 77.8437795956, 26.8299799704, 35.0000346037, 35.9651027691};
test_label[2235] = '{35.9651027691};
test_output[2235] = '{57.9292000986};
############ END DEBUG ############*/
test_input[17888:17895] = '{32'h416cfa3e, 32'hc275eac9, 32'h42aea3e4, 32'hc26a25bf, 32'h42888940, 32'hc226e7b3, 32'h42c0060a, 32'hc10b1589};
test_label[2236] = '{32'hc226e7b3};
test_output[2236] = '{32'h4309bcfd};
/*############ DEBUG ############
test_input[17888:17895] = '{14.8110940947, -61.4792825487, 87.3200990199, -58.5368613404, 68.2680684001, -41.7262698526, 96.0117914046, -8.69275743758};
test_label[2236] = '{-41.7262698526};
test_output[2236] = '{137.738229219};
############ END DEBUG ############*/
test_input[17896:17903] = '{32'h42b2875c, 32'hc1f66153, 32'hc1952396, 32'h42173ad6, 32'hc1891c6b, 32'h42c6d53d, 32'h426894e2, 32'h412aa87d};
test_label[2237] = '{32'hc1891c6b};
test_output[2237] = '{32'h42e91c5d};
/*############ DEBUG ############
test_input[17896:17903] = '{89.2643711551, -30.797521897, -18.6423756725, 37.8074567502, -17.1388755146, 99.4164833243, 58.1453949092, 10.6661350677};
test_label[2237] = '{-17.1388755146};
test_output[2237] = '{116.555397832};
############ END DEBUG ############*/
test_input[17904:17911] = '{32'hc22af999, 32'h4210a25a, 32'hc2c334bd, 32'h4208ac49, 32'h42b53a72, 32'hc28ee8ae, 32'hc2c2a5a7, 32'h422dd7c8};
test_label[2238] = '{32'hc2c334bd};
test_output[2238] = '{32'h433c3798};
/*############ DEBUG ############
test_input[17904:17911] = '{-42.7437494123, 36.1585451421, -97.603005949, 34.1682474727, 90.614153691, -71.4544497856, -97.3235388078, 43.4607225858};
test_label[2238] = '{-97.603005949};
test_output[2238] = '{188.21715964};
############ END DEBUG ############*/
test_input[17912:17919] = '{32'h41fe3517, 32'h422bbced, 32'h42b20616, 32'hc2b4ea5f, 32'h42248e36, 32'hc245ffa1, 32'h3f5dec8d, 32'hc298325a};
test_label[2239] = '{32'h422bbced};
test_output[2239] = '{32'h42384f3e};
/*############ DEBUG ############
test_input[17912:17919] = '{31.7759232284, 42.9344974903, 89.0118829726, -90.457752555, 41.1388772557, -49.4996379817, 0.866890740884, -76.0983400223};
test_label[2239] = '{42.9344974903};
test_output[2239] = '{46.0773854824};
############ END DEBUG ############*/
test_input[17920:17927] = '{32'h429a185f, 32'h411453f3, 32'hc21ebd4b, 32'hc2b0aedf, 32'hc1ada3a8, 32'hc183ce3e, 32'h4292ff6f, 32'h3eb1fee5};
test_label[2240] = '{32'hc21ebd4b};
test_output[2240] = '{32'h42e98589};
/*############ DEBUG ############
test_input[17920:17927] = '{77.0475964004, 9.27049559671, -39.6848553526, -88.3415413932, -21.7049104901, -16.4757048333, 73.4988905679, 0.347647807176};
test_label[2240] = '{-39.6848553526};
test_output[2240] = '{116.760807733};
############ END DEBUG ############*/
test_input[17928:17935] = '{32'h42833148, 32'h428d6f3a, 32'h4166bb3e, 32'hc286e47b, 32'h42aaac51, 32'hc2188676, 32'h4284d2f7, 32'h41fc175a};
test_label[2241] = '{32'hc2188676};
test_output[2241] = '{32'h42f6ef8c};
/*############ DEBUG ############
test_input[17928:17935] = '{65.5962523265, 70.7172429257, 14.4207132456, -67.4462501944, 85.3365531744, -38.1313109443, 66.4120391294, 31.5114024683};
test_label[2241] = '{-38.1313109443};
test_output[2241] = '{123.467864575};
############ END DEBUG ############*/
test_input[17936:17943] = '{32'hc22c78e6, 32'h41b6bb41, 32'h428328a7, 32'h424787c2, 32'h410e00c5, 32'hc27a3332, 32'hc127571b, 32'hc1d58b0a};
test_label[2242] = '{32'hc27a3332};
test_output[2242] = '{32'h43002120};
/*############ DEBUG ############
test_input[17936:17943] = '{-43.118066193, 22.841431752, 65.5793962625, 49.8825747459, 8.87518780536, -62.5499950746, -10.4587656276, -26.6928900221};
test_label[2242] = '{-62.5499950746};
test_output[2242] = '{128.12939149};
############ END DEBUG ############*/
test_input[17944:17951] = '{32'h4229dac3, 32'hc21b6da5, 32'h40e047b7, 32'hc215981c, 32'h42a54a5f, 32'hc2164037, 32'hc2be3568, 32'hc1ffdfcf};
test_label[2243] = '{32'hc21b6da5};
test_output[2243] = '{32'h42f30132};
/*############ DEBUG ############
test_input[17944:17951] = '{42.4636342704, -38.8570765396, 7.00875434716, -37.3985424929, 82.6452547287, -37.5627088336, -95.1043109752, -31.9842807396};
test_label[2243] = '{-38.8570765396};
test_output[2243] = '{121.502331268};
############ END DEBUG ############*/
test_input[17952:17959] = '{32'hc2a35a6e, 32'h421b52cf, 32'hc26d188f, 32'h418d868f, 32'h422deb6c, 32'hc23eaea4, 32'h41b5b44a, 32'h42060058};
test_label[2244] = '{32'h41b5b44a};
test_output[2244] = '{32'h41a63628};
/*############ DEBUG ############
test_input[17952:17959] = '{-81.6766234526, 38.8308672191, -59.2739839716, 17.6907029828, 43.4799047503, -47.6705466061, 22.713032286, 33.5003350158};
test_label[2244] = '{22.713032286};
test_output[2244] = '{20.776443661};
############ END DEBUG ############*/
test_input[17960:17967] = '{32'h429fccb8, 32'h4253b31f, 32'hc293f264, 32'h42c067ef, 32'hc2b19360, 32'h426f8440, 32'h42b74135, 32'hc29a6a49};
test_label[2245] = '{32'h426f8440};
test_output[2245] = '{32'h4211561d};
/*############ DEBUG ############
test_input[17960:17967] = '{79.8998400732, 52.9249211564, -73.9734183878, 96.2029965176, -88.7878393633, 59.879149186, 91.6273548983, -77.2075861141};
test_label[2245] = '{59.879149186};
test_output[2245] = '{36.3340944221};
############ END DEBUG ############*/
test_input[17968:17975] = '{32'hc2c26ae6, 32'hc2ac2cb8, 32'h42b6d7f0, 32'hc2a73765, 32'hc2c6e23b, 32'hc1b5f87d, 32'hc2978fa7, 32'h419a43dc};
test_label[2246] = '{32'hc2c26ae6};
test_output[2246] = '{32'h433ca16b};
/*############ DEBUG ############
test_input[17968:17975] = '{-97.2087847347, -86.0873442593, 91.4217530619, -83.6081949008, -99.4418548439, -22.7463328913, -75.7805716296, 19.2831348779};
test_label[2246] = '{-97.2087847347};
test_output[2246] = '{188.630537797};
############ END DEBUG ############*/
test_input[17976:17983] = '{32'hc27d76f2, 32'h4000570f, 32'hc21f174c, 32'h429ec47b, 32'h42a78e77, 32'h42bd6b92, 32'hc1e901dc, 32'hc2405c19};
test_label[2247] = '{32'hc2405c19};
test_output[2247] = '{32'h430eccd0};
/*############ DEBUG ############
test_input[17976:17983] = '{-63.3661571078, 2.00531369664, -39.772749014, 79.3837526467, 83.7782532183, 94.7100967983, -29.1259087401, -48.0899383953};
test_label[2247] = '{-48.0899383953};
test_output[2247] = '{142.800053294};
############ END DEBUG ############*/
test_input[17984:17991] = '{32'hc15ba9e9, 32'h413e0059, 32'hc1b79606, 32'hc1b19b27, 32'h4251985b, 32'h420a4eff, 32'h425a3933, 32'h406650d4};
test_label[2248] = '{32'h406650d4};
test_output[2248] = '{32'h424c4439};
/*############ DEBUG ############
test_input[17984:17991] = '{-13.7289816613, 11.8750851924, -22.9482534584, -22.2007585849, 52.3987841852, 34.5771438621, 54.5558586485, 3.59868338541};
test_label[2248] = '{3.59868338541};
test_output[2248] = '{51.0666241146};
############ END DEBUG ############*/
test_input[17992:17999] = '{32'hc20507d6, 32'hc29c0de1, 32'hc2291095, 32'hc23c6d75, 32'hc2159abf, 32'h424866f2, 32'hc2acd3ab, 32'h42a1d0c6};
test_label[2249] = '{32'hc23c6d75};
test_output[2249] = '{32'h430003c0};
/*############ DEBUG ############
test_input[17992:17999] = '{-33.2576534746, -78.0271064268, -42.266191892, -47.1068898885, -37.4011184448, 50.100532122, -86.4134144767, 80.9077584175};
test_label[2249] = '{-47.1068898885};
test_output[2249] = '{128.014648306};
############ END DEBUG ############*/
test_input[18000:18007] = '{32'hc2b8518f, 32'hc2086349, 32'h428ebe61, 32'hc24c36b4, 32'h42c76588, 32'h42587b9a, 32'hc25bbf8a, 32'h41c918e7};
test_label[2250] = '{32'hc2b8518f};
test_output[2250] = '{32'h433fdb8b};
/*############ DEBUG ############
test_input[18000:18007] = '{-92.1592935862, -34.0969572083, 71.3718330311, -51.0534202926, 99.6983010753, 54.1207034383, -54.937048188, 25.1371601476};
test_label[2250] = '{-92.1592935862};
test_output[2250] = '{191.857594661};
############ END DEBUG ############*/
test_input[18008:18015] = '{32'h4271b8c5, 32'hc2360714, 32'h404c6efa, 32'hc2a88c1a, 32'h41854952, 32'hc2872064, 32'hc2b569bf, 32'hc262cea2};
test_label[2251] = '{32'hc262cea2};
test_output[2251] = '{32'h42ea43b4};
/*############ DEBUG ############
test_input[18008:18015] = '{60.4304407032, -45.5069131251, 3.19427339614, -84.2736332633, 16.660801844, -67.563265436, -90.7065342668, -56.7017886856};
test_label[2251] = '{-56.7017886856};
test_output[2251] = '{117.132229389};
############ END DEBUG ############*/
test_input[18016:18023] = '{32'h42934121, 32'h42469cdf, 32'h4115144e, 32'hc2482e39, 32'hc1484f61, 32'h425667ba, 32'hc1292541, 32'hc2b33fc3};
test_label[2252] = '{32'h42934121};
test_output[2252] = '{32'h310cae76};
/*############ DEBUG ############
test_input[18016:18023] = '{73.6272027881, 49.6531942077, 9.31745752707, -50.0451376965, -12.5193793237, 53.6012951377, -10.5715949498, -89.624533687};
test_label[2252] = '{73.6272027881};
test_output[2252] = '{2.04718509021e-09};
############ END DEBUG ############*/
test_input[18024:18031] = '{32'h4262fccb, 32'h4240e147, 32'h421c5f70, 32'h42905485, 32'h41fc2ed5, 32'hc1e35016, 32'h4287109e, 32'hc2a9cc82};
test_label[2253] = '{32'h4262fccb};
test_output[2253] = '{32'h4176d8a4};
/*############ DEBUG ############
test_input[18024:18031] = '{56.7468696235, 48.2199978487, 39.0932024867, 72.1650782876, 31.5228665995, -28.4141040796, 67.5324549334, -84.8994295481};
test_label[2253] = '{56.7468696235};
test_output[2253] = '{15.4278910421};
############ END DEBUG ############*/
test_input[18032:18039] = '{32'hc2079af8, 32'hc28bbb32, 32'h41ae0271, 32'h42b4ce77, 32'hc22061df, 32'hc2b40476, 32'hc2285e76, 32'hc2ba6f07};
test_label[2254] = '{32'hc28bbb32};
test_output[2254] = '{32'h432044d4};
/*############ DEBUG ############
test_input[18032:18039] = '{-33.9013380891, -69.8656143246, 21.7511916637, 90.4032481098, -40.0955755222, -90.0087151904, -42.0922488204, -93.2168512842};
test_label[2254] = '{-69.8656143246};
test_output[2254] = '{160.268862434};
############ END DEBUG ############*/
test_input[18040:18047] = '{32'h40b33caa, 32'hc285e168, 32'hc2554cde, 32'hc1cb1e9b, 32'h42005b63, 32'h42ba8e87, 32'hc2bc6b4c, 32'h4294b355};
test_label[2255] = '{32'h42ba8e87};
test_output[2255] = '{32'h31cedbcc};
/*############ DEBUG ############
test_input[18040:18047] = '{5.60115510087, -66.9402447712, -53.3250646535, -25.3899442342, 32.0892437937, 93.2783768556, -94.2095630152, 74.350260926};
test_label[2255] = '{93.2783768556};
test_output[2255] = '{6.02037710387e-09};
############ END DEBUG ############*/
test_input[18048:18055] = '{32'hc29e41c7, 32'hbfac59fe, 32'hc1fb7d47, 32'hc23d1751, 32'h41dc7f90, 32'hc26586bc, 32'h4212f4db, 32'h42a3b96d};
test_label[2256] = '{32'h4212f4db};
test_output[2256] = '{32'h42347dff};
/*############ DEBUG ############
test_input[18048:18055] = '{-79.1284740291, -1.34649629017, -31.4361706834, -47.2727692066, 27.5622868374, -57.3815766234, 36.739117295, 81.8621603499};
test_label[2256] = '{36.739117295};
test_output[2256] = '{45.1230430549};
############ END DEBUG ############*/
test_input[18056:18063] = '{32'hc2b083f8, 32'hc2856e33, 32'hc1d40c4a, 32'hc26c15a6, 32'h422ead9c, 32'h41fc1262, 32'hc29a61f1, 32'hc27814fb};
test_label[2257] = '{32'h41fc1262};
test_output[2257] = '{32'h414291b1};
/*############ DEBUG ############
test_input[18056:18063] = '{-88.2577477655, -66.7152302012, -26.5059998747, -59.0211409712, 43.6695391478, 31.5089751412, -77.1912918354, -62.0204876968};
test_label[2257] = '{31.5089751412};
test_output[2257] = '{12.1605692394};
############ END DEBUG ############*/
test_input[18064:18071] = '{32'hc2253472, 32'h42a1ace6, 32'hc2c4004f, 32'h4197fda3, 32'h41be3b5f, 32'hc2c45474, 32'h41cae7de, 32'hc1f1aba6};
test_label[2258] = '{32'hc1f1aba6};
test_output[2258] = '{32'h42de17d0};
/*############ DEBUG ############
test_input[18064:18071] = '{-41.3012171896, 80.8376957602, -98.0006027622, 18.9988464296, 23.7789891762, -98.164946831, 25.3632169582, -30.2088124267};
test_label[2258] = '{-30.2088124267};
test_output[2258] = '{111.046508187};
############ END DEBUG ############*/
test_input[18072:18079] = '{32'hc289bbd9, 32'h426ba093, 32'h42845e2c, 32'h423bfe7c, 32'h42b471fd, 32'hc152bd4d, 32'h42a52ef4, 32'h429e1134};
test_label[2259] = '{32'h426ba093};
test_output[2259] = '{32'h41fa87d3};
/*############ DEBUG ############
test_input[18072:18079] = '{-68.866891735, 58.9068095574, 66.1839319271, 46.9985207735, 90.2226311278, -13.1712157514, 82.5917043278, 79.0335995326};
test_label[2259] = '{58.9068095574};
test_output[2259] = '{31.316320482};
############ END DEBUG ############*/
test_input[18080:18087] = '{32'h42c4150f, 32'hc29d44b9, 32'hc289c1e1, 32'hc23fbc97, 32'h423353fd, 32'h427d4d93, 32'h42c3724d, 32'hc2235643};
test_label[2260] = '{32'hc29d44b9};
test_output[2260] = '{32'h433138de};
/*############ DEBUG ############
test_input[18080:18087] = '{98.0411289259, -78.6342259729, -68.8786711515, -47.9341687893, 44.832019019, 63.3257546155, 97.7232423603, -40.8342381189};
test_label[2260] = '{-78.6342259729};
test_output[2260] = '{177.222137451};
############ END DEBUG ############*/
test_input[18088:18095] = '{32'hc2bb2b40, 32'hc1e6d046, 32'hc2c64d67, 32'hc1d26f37, 32'hc15f8269, 32'h41c3a778, 32'hc29c0e00, 32'h429b06a9};
test_label[2261] = '{32'h429b06a9};
test_output[2261] = '{32'h80000000};
/*############ DEBUG ############
test_input[18088:18095] = '{-93.5844751274, -28.8516951624, -99.1511767196, -26.3043050249, -13.9693380685, 24.4567711115, -78.0273429235, 77.5130081478};
test_label[2261] = '{77.5130081478};
test_output[2261] = '{-0.0};
############ END DEBUG ############*/
test_input[18096:18103] = '{32'hc22f8a22, 32'h42bc9190, 32'h42acdc71, 32'hc220bd31, 32'h42220a58, 32'hc2992064, 32'hc2bb5d27, 32'hc1b0d0b0};
test_label[2262] = '{32'hc1b0d0b0};
test_output[2262] = '{32'h42e8c5ef};
/*############ DEBUG ############
test_input[18096:18103] = '{-43.8848953764, 94.284304551, 86.4305463292, -40.1847571983, 40.5100997832, -76.5632593887, -93.6819353608, -22.1018982716};
test_label[2262] = '{-22.1018982716};
test_output[2262] = '{116.386591037};
############ END DEBUG ############*/
test_input[18104:18111] = '{32'h4269a3ae, 32'h420c94ff, 32'hc19f6f35, 32'h42329461, 32'hc1b809c0, 32'h429efcf0, 32'hc28e6d4f, 32'hc1447d8e};
test_label[2263] = '{32'hc19f6f35};
test_output[2263] = '{32'h42c6d8bd};
/*############ DEBUG ############
test_input[18104:18111] = '{58.4098428354, 35.1455021304, -19.9293004854, 44.6449027898, -23.0047604716, 79.4940179421, -71.2134949628, -12.280652578};
test_label[2263] = '{-19.9293004854};
test_output[2263] = '{99.4233184282};
############ END DEBUG ############*/
test_input[18112:18119] = '{32'h418bd215, 32'hc29c3458, 32'hc298ea2c, 32'hc20c3342, 32'hc2263990, 32'h42a1310b, 32'hc1e13236, 32'h41b8dd35};
test_label[2264] = '{32'hc2263990};
test_output[2264] = '{32'h42f44dd3};
/*############ DEBUG ############
test_input[18112:18119] = '{17.4775799278, -78.1022307319, -76.4573684803, -35.0500570118, -41.556214638, 80.5957895776, -28.149517137, 23.1080121542};
test_label[2264] = '{-41.556214638};
test_output[2264] = '{122.152004216};
############ END DEBUG ############*/
test_input[18120:18127] = '{32'h42467236, 32'h4297157d, 32'h420455db, 32'hc287c33f, 32'h426e3980, 32'h42b2a201, 32'h421773bc, 32'hc2b398c5};
test_label[2265] = '{32'h42b2a201};
test_output[2265] = '{32'h358bd826};
/*############ DEBUG ############
test_input[18120:18127] = '{49.6115340702, 75.5419672967, 33.0838429039, -67.8813380389, 59.5561513461, 89.3164108449, 37.8630218335, -89.7983781371};
test_label[2265] = '{89.3164108449};
test_output[2265] = '{1.04192149831e-06};
############ END DEBUG ############*/
test_input[18128:18135] = '{32'h4264800c, 32'hc2a26b3a, 32'h42264bd8, 32'hc2a3c99f, 32'hc28de3b3, 32'h427ecc66, 32'hc2b6a49a, 32'h401feb83};
test_label[2266] = '{32'h42264bd8};
test_output[2266] = '{32'h41b103f8};
/*############ DEBUG ############
test_input[18128:18135] = '{57.1250451992, -81.2094287151, 41.5740646108, -81.8937906956, -70.9447217754, 63.6996073568, -91.3214850088, 2.49874953604};
test_label[2266] = '{41.5740646108};
test_output[2266] = '{22.1269371903};
############ END DEBUG ############*/
test_input[18136:18143] = '{32'h420f1cbb, 32'h42bb0b2c, 32'h41a94283, 32'h42b5229d, 32'hc0f84cc4, 32'h4287e6b0, 32'hc2c68b9e, 32'hc284b1f5};
test_label[2267] = '{32'h4287e6b0};
test_output[2267] = '{32'h41ccf9fc};
/*############ DEBUG ############
test_input[18136:18143] = '{35.7780583663, 93.5218192445, 21.1574759554, 90.5676051222, -7.75937070845, 67.9505639292, -99.2726927483, -66.3475691941};
test_label[2267] = '{67.9505639292};
test_output[2267] = '{25.6220621153};
############ END DEBUG ############*/
test_input[18144:18151] = '{32'hc2bfc815, 32'h41c0f360, 32'h428901fb, 32'h4223d6bd, 32'h411d96b3, 32'h429a6861, 32'h4163c649, 32'h42b4ec54};
test_label[2268] = '{32'hc2bfc815};
test_output[2268] = '{32'h433a5a34};
/*############ DEBUG ############
test_input[18144:18151] = '{-95.8907830944, 24.1188355494, 68.5038667893, 40.9597043447, 9.84929136976, 77.2038687081, 14.2359090164, 90.461577167};
test_label[2268] = '{-95.8907830944};
test_output[2268] = '{186.352362009};
############ END DEBUG ############*/
test_input[18152:18159] = '{32'hc219e04d, 32'h4291c30d, 32'hc2902c0b, 32'hc273eaa6, 32'hc29abd95, 32'hc249e213, 32'h42a8aaea, 32'hbd94312b};
test_label[2269] = '{32'h4291c30d};
test_output[2269] = '{32'h41373ef5};
/*############ DEBUG ############
test_input[18152:18159] = '{-38.4690424564, 72.8809561457, -72.0860192807, -60.9791488808, -77.3702740677, -50.4707751037, 84.3338156684, -0.0723594077581};
test_label[2269] = '{72.8809561457};
test_output[2269] = '{11.4528701417};
############ END DEBUG ############*/
test_input[18160:18167] = '{32'h426ac61e, 32'hc129f54f, 32'h41fdf83b, 32'h4277cb22, 32'hc293ee1c, 32'hc2badad0, 32'h42b04b8b, 32'h42c7b016};
test_label[2270] = '{32'hc293ee1c};
test_output[2270] = '{32'h432dcf1a};
/*############ DEBUG ############
test_input[18160:18167] = '{58.6934724374, -10.6223897428, 31.7462055185, 61.9483727254, -73.9650560697, -93.427369826, 88.1475478186, 99.8439186364};
test_label[2270] = '{-73.9650560697};
test_output[2270] = '{173.80898303};
############ END DEBUG ############*/
test_input[18168:18175] = '{32'hc189d66d, 32'h41764293, 32'hc1a8abcb, 32'h41c48d59, 32'hc2320305, 32'hc24ffdd3, 32'h41a94565, 32'hc29f0467};
test_label[2271] = '{32'hc24ffdd3};
test_output[2271] = '{32'h429932f1};
/*############ DEBUG ############
test_input[18168:18175] = '{-17.2296993631, 15.3912530779, -21.083883046, 24.5690166093, -44.5029505437, -51.997875442, 21.1588831719, -79.5085989165};
test_label[2271] = '{-51.997875442};
test_output[2271] = '{76.5994948595};
############ END DEBUG ############*/
test_input[18176:18183] = '{32'hc267eba5, 32'h425f0c39, 32'h411f9082, 32'h42a39901, 32'hc26bd46f, 32'hc02b553a, 32'hc25442a0, 32'h41abccd2};
test_label[2272] = '{32'hc26bd46f};
test_output[2272] = '{32'h430cc19d};
/*############ DEBUG ############
test_input[18176:18183] = '{-57.9801203195, 55.7619379326, 9.97278064142, 81.7988393327, -58.9574563317, -2.67707683927, -53.0650645429, 21.4750090244};
test_label[2272] = '{-58.9574563317};
test_output[2272] = '{140.756295664};
############ END DEBUG ############*/
test_input[18184:18191] = '{32'hc256c37c, 32'hc2148546, 32'hc2b64eda, 32'h429ea098, 32'h425ff585, 32'hc1081e8d, 32'hc19084c3, 32'hc1f1d0c3};
test_label[2273] = '{32'hc19084c3};
test_output[2273] = '{32'h42c2c1c9};
/*############ DEBUG ############
test_input[18184:18191] = '{-53.6909042384, -37.130147983, -91.1540049537, 79.313659563, 55.9897655023, -8.50745887156, -18.0648255599, -30.2269347867};
test_label[2273] = '{-18.0648255599};
test_output[2273] = '{97.378485123};
############ END DEBUG ############*/
test_input[18192:18199] = '{32'h4192d6eb, 32'hc18090e1, 32'hc2be9e54, 32'hc2480579, 32'hc147802f, 32'h42c573ec, 32'hc2c7b9fd, 32'hc28f45d6};
test_label[2274] = '{32'hc2c7b9fd};
test_output[2274] = '{32'h434696f4};
/*############ DEBUG ############
test_input[18192:18199] = '{18.3549409966, -16.0707419002, -95.3092361362, -50.0053459043, -12.4687948637, 98.7264101665, -99.8632569325, -71.6364005288};
test_label[2274] = '{-99.8632569325};
test_output[2274] = '{198.589667099};
############ END DEBUG ############*/
test_input[18200:18207] = '{32'h4295138b, 32'h4282c664, 32'hc2883725, 32'h42665bd6, 32'hc194e352, 32'hc22285bc, 32'hc1849284, 32'h427a4041};
test_label[2275] = '{32'hc194e352};
test_output[2275] = '{32'h42ba4c6f};
/*############ DEBUG ############
test_input[18200:18207] = '{74.5381733486, 65.3874848332, -68.1077066125, 57.5896846658, -18.6109962927, -40.6305982751, -16.5715415107, 62.562747239};
test_label[2275] = '{-18.6109962927};
test_output[2275] = '{93.1492821224};
############ END DEBUG ############*/
test_input[18208:18215] = '{32'h41d9e01e, 32'h417ec9ef, 32'hc2b0bb7e, 32'h426751d3, 32'h42bda784, 32'h420bf69c, 32'h419a480f, 32'h41079dcc};
test_label[2276] = '{32'h426751d3};
test_output[2276] = '{32'h4213fd35};
/*############ DEBUG ############
test_input[18208:18215] = '{27.2344320811, 15.9243002681, -88.366197134, 57.8299074684, 94.8271790042, 34.9908295944, 19.2851841775, 8.47602486146};
test_label[2276] = '{57.8299074684};
test_output[2276] = '{36.9972715358};
############ END DEBUG ############*/
test_input[18216:18223] = '{32'h423252de, 32'h41cf74ba, 32'hc29c3f3d, 32'hc0081e7b, 32'hc2bc6b26, 32'h4271efb2, 32'h429c2ead, 32'h4171a4cf};
test_label[2277] = '{32'h4271efb2};
test_output[2277] = '{32'h418cdb4e};
/*############ DEBUG ############
test_input[18216:18223] = '{44.5809253015, 25.9319955187, -78.1235106461, -2.12686035015, -94.2092721864, 60.4840778462, 78.0911604, 15.1027364088};
test_label[2277] = '{60.4840778462};
test_output[2277] = '{17.6070825763};
############ END DEBUG ############*/
test_input[18224:18231] = '{32'hc22a67b0, 32'h429e5380, 32'h42942297, 32'hc2937ce9, 32'hc289ffb9, 32'h42a2fdfd, 32'hc2786179, 32'hc2a64b16};
test_label[2278] = '{32'hc2a64b16};
test_output[2278] = '{32'h4324bc61};
/*############ DEBUG ############
test_input[18224:18231] = '{-42.6012589911, 79.163087013, 74.0675560113, -73.7439668551, -68.9994568702, 81.4960734954, -62.095188667, -83.1466544124};
test_label[2278] = '{-83.1466544124};
test_output[2278] = '{164.735853591};
############ END DEBUG ############*/
test_input[18232:18239] = '{32'hc1b6a7d7, 32'hc2731cdf, 32'h42b36b9a, 32'h42a9f789, 32'h4292beb3, 32'h4289a3ef, 32'h422b84e6, 32'hc145d103};
test_label[2279] = '{32'hc1b6a7d7};
test_output[2279] = '{32'h42e11a13};
/*############ DEBUG ############
test_input[18232:18239] = '{-22.831952109, -60.7781927046, 89.7101595358, 84.9834675574, 73.3724569035, 68.8201839596, 42.8797819531, -12.363528717};
test_label[2279] = '{-22.831952109};
test_output[2279] = '{112.550928461};
############ END DEBUG ############*/
test_input[18240:18247] = '{32'h429aac21, 32'h426c9d7d, 32'h42ba3d4f, 32'hc2306b7b, 32'h40b5a9bd, 32'h420dabcb, 32'hc134afdf, 32'hc1ec9e23};
test_label[2280] = '{32'hc2306b7b};
test_output[2280] = '{32'h43093987};
/*############ DEBUG ############
test_input[18240:18247] = '{77.3361923375, 59.1537960437, 93.1197465358, -44.1049626055, 5.67697019037, 35.4177651217, -11.2929373132, -29.5772145708};
test_label[2280] = '{-44.1049626055};
test_output[2280] = '{137.224709281};
############ END DEBUG ############*/
test_input[18248:18255] = '{32'hc2847871, 32'hc2b68f00, 32'h419fe3dc, 32'hc2642f53, 32'h4291a4f6, 32'h40714096, 32'hc1c89b18, 32'h4213d85d};
test_label[2281] = '{32'h4213d85d};
test_output[2281] = '{32'h420f718e};
/*############ DEBUG ############
test_input[18248:18255] = '{-66.2352362642, -91.2792943058, 19.9862602434, -57.0462152704, 72.8221863912, 3.76956701095, -25.075728659, 36.9612933775};
test_label[2281] = '{36.9612933775};
test_output[2281] = '{35.8608930136};
############ END DEBUG ############*/
test_input[18256:18263] = '{32'hc2b0e5be, 32'hc2b2f86c, 32'h4280f8d3, 32'h4174d98e, 32'hc2b6302c, 32'h42c287d6, 32'h428ef488, 32'h41a34fbf};
test_label[2282] = '{32'hc2b2f86c};
test_output[2282] = '{32'h433ac021};
/*############ DEBUG ############
test_input[18256:18263] = '{-88.4487166018, -89.4852006457, 64.4859835778, 15.30311362, -91.0940893663, 97.2653045562, 71.4776011012, 20.4139384152};
test_label[2282] = '{-89.4852006457};
test_output[2282] = '{186.750505202};
############ END DEBUG ############*/
test_input[18264:18271] = '{32'hc14209e9, 32'hc28ddc82, 32'h42807320, 32'h4288b200, 32'hc2a9edaa, 32'h3fdcdd3c, 32'h429b609d, 32'hc2c064f6};
test_label[2283] = '{32'h3fdcdd3c};
test_output[2283] = '{32'h4297ed33};
/*############ DEBUG ############
test_input[18264:18271] = '{-12.1274195212, -70.9306814024, 64.2248569718, 68.3476570179, -84.9641909603, 1.72550151901, 77.6886948649, -96.1971879329};
test_label[2283] = '{1.72550151901};
test_output[2283] = '{75.9632825117};
############ END DEBUG ############*/
test_input[18272:18279] = '{32'h4235163c, 32'h4183dbf1, 32'h411b93bb, 32'hc2930658, 32'h41a1caae, 32'h423e3389, 32'h4239d1d7, 32'h3f998ce2};
test_label[2284] = '{32'h4239d1d7};
test_output[2284] = '{32'h3fba9aa0};
/*############ DEBUG ############
test_input[18272:18279] = '{45.2717131491, 16.4823933576, 9.72356740992, -73.5123868871, 20.2239654754, 47.5503264692, 46.454922447, 1.19961187172};
test_label[2284] = '{46.454922447};
test_output[2284] = '{1.45784374717};
############ END DEBUG ############*/
test_input[18280:18287] = '{32'h420d4c0c, 32'hc2bf2db9, 32'hbdc2205e, 32'h4283befb, 32'hc21648dd, 32'hc1f8ad63, 32'h414b4046, 32'hc293b615};
test_label[2285] = '{32'hc1f8ad63};
test_output[2285] = '{32'h42c1ea53};
/*############ DEBUG ############
test_input[18280:18287] = '{35.3242648111, -95.5893048339, -0.0947882993584, 65.8730055826, -37.5711561808, -31.0846605778, 12.7031922201, -73.855626729};
test_label[2285] = '{-31.0846605778};
test_output[2285] = '{96.9576661604};
############ END DEBUG ############*/
test_input[18288:18295] = '{32'h4288213f, 32'h427f608c, 32'hc1124e9c, 32'h42c72d36, 32'h4286d64b, 32'hc2aa9e0b, 32'hc2887c72, 32'h42aabfa5};
test_label[2286] = '{32'h4286d64b};
test_output[2286] = '{32'h4200add6};
/*############ DEBUG ############
test_input[18288:18295] = '{68.0649322798, 63.8442845316, -9.14419147558, 99.5882996845, 67.4185371469, -85.3086796807, -68.2430543765, 85.3743052645};
test_label[2286] = '{67.4185371469};
test_output[2286] = '{32.1697632089};
############ END DEBUG ############*/
test_input[18296:18303] = '{32'h42a3b468, 32'h42c44eb2, 32'hc24183df, 32'hc2bc6c67, 32'hc2a9f576, 32'hc2b5231b, 32'h422ec0d1, 32'hc2994727};
test_label[2287] = '{32'h42c44eb2};
test_output[2287] = '{32'h33b2ca46};
/*############ DEBUG ############
test_input[18296:18303] = '{81.8523540628, 98.1537039734, -48.3787808781, -94.2117270537, -84.9794142704, -90.5685625085, 43.688298317, -76.6389717729};
test_label[2287] = '{98.1537039734};
test_output[2287] = '{8.325564085e-08};
############ END DEBUG ############*/
test_input[18304:18311] = '{32'h4292c875, 32'hc1076cf5, 32'hc01e028c, 32'hc2b125a5, 32'h42956690, 32'h41fea957, 32'h42a815a2, 32'hc294e0b8};
test_label[2288] = '{32'h42956690};
test_output[2288] = '{32'h41157901};
/*############ DEBUG ############
test_input[18304:18311] = '{73.3915151453, -8.46410108251, -2.4689054828, -88.5735229619, 74.7003189253, 31.8326856848, 84.0422491326, -74.4389047427};
test_label[2288] = '{74.7003189253};
test_output[2288] = '{9.34204155464};
############ END DEBUG ############*/
test_input[18312:18319] = '{32'hc251eec8, 32'h428c0895, 32'h420c881c, 32'hc22e416e, 32'hc29052b4, 32'hc2b25540, 32'h40a0750f, 32'hc248e4e7};
test_label[2289] = '{32'hc22e416e};
test_output[2289] = '{32'h42e3294c};
/*############ DEBUG ############
test_input[18312:18319] = '{-52.4831829322, 70.0167650451, 35.1329193836, -43.5638945209, -72.1615290964, -89.1665053035, 5.01428929754, -50.2235384235};
test_label[2289] = '{-43.5638945209};
test_output[2289] = '{113.580659566};
############ END DEBUG ############*/
test_input[18320:18327] = '{32'hc1cb232c, 32'h42a23752, 32'h42968a80, 32'h428f2aa4, 32'hc1a869d4, 32'hc12e1aeb, 32'hc19a0f07, 32'hc278eb48};
test_label[2290] = '{32'hc1cb232c};
test_output[2290] = '{32'h42d501a4};
/*############ DEBUG ############
test_input[18320:18327] = '{-25.3921731424, 81.1080471202, 75.270506866, 71.5832829634, -21.0516745605, -10.8815714214, -19.2573379657, -62.2297655151};
test_label[2290] = '{-25.3921731424};
test_output[2290] = '{106.503204832};
############ END DEBUG ############*/
test_input[18328:18335] = '{32'h42b11b76, 32'h4289026a, 32'h410a713b, 32'h421e26da, 32'hc2a7e074, 32'h4102b6c7, 32'h425f11fe, 32'h42931cc1};
test_label[2291] = '{32'hc2a7e074};
test_output[2291] = '{32'h432c7df5};
/*############ DEBUG ############
test_input[18328:18335] = '{88.5536364604, 68.5047168563, 8.65264441452, 39.5379427968, -83.9383869402, 8.16962324624, 55.7675714339, 73.5561610955};
test_label[2291] = '{-83.9383869402};
test_output[2291] = '{172.492023709};
############ END DEBUG ############*/
test_input[18336:18343] = '{32'hc1de70ee, 32'hc2bfc71d, 32'h4191c621, 32'h4268d67e, 32'hc286f0be, 32'hc24c5f15, 32'hc21511f1, 32'h42bde5e5};
test_label[2292] = '{32'hc21511f1};
test_output[2292] = '{32'h4304376f};
/*############ DEBUG ############
test_input[18336:18343] = '{-27.8051413838, -95.8888925827, 18.2217429581, 58.2094634948, -67.4702015089, -51.0928531474, -37.2675209193, 94.9490128756};
test_label[2292] = '{-37.2675209193};
test_output[2292] = '{132.216533795};
############ END DEBUG ############*/
test_input[18344:18351] = '{32'h41babb9f, 32'hc297cc94, 32'hc258d258, 32'h41b47526, 32'hc2849efd, 32'h410651a6, 32'h42b240c3, 32'h42bfe399};
test_label[2293] = '{32'h42bfe399};
test_output[2293] = '{32'h3a8f4bf7};
/*############ DEBUG ############
test_input[18344:18351] = '{23.3416116633, -75.8995631274, -54.2054131958, 22.557201021, -66.3105228782, 8.39493341023, 89.1264906754, 95.9445285043};
test_label[2293] = '{95.9445285043};
test_output[2293] = '{0.00109326733394};
############ END DEBUG ############*/
test_input[18352:18359] = '{32'h41cbec2e, 32'h41061ef0, 32'h429205c1, 32'hc2181fa4, 32'h415a9bba, 32'hc26bb91e, 32'h41afa400, 32'h41ec56ec};
test_label[2294] = '{32'h41061ef0};
test_output[2294] = '{32'h428141e3};
/*############ DEBUG ############
test_input[18352:18359] = '{25.4903220978, 8.38255345301, 73.0112396009, -38.0308983715, 13.6630194968, -58.9307769636, 21.9550775221, 29.5424426453};
test_label[2294] = '{8.38255345301};
test_output[2294] = '{64.6286861479};
############ END DEBUG ############*/
test_input[18360:18367] = '{32'h42ae735f, 32'hc28ee6c6, 32'hc298d8e7, 32'h41e64177, 32'h42a74cd7, 32'h42775bab, 32'h4278701e, 32'hc1df6f09};
test_label[2295] = '{32'h42ae735f};
test_output[2295] = '{32'h3ce249dd};
/*############ DEBUG ############
test_input[18360:18367] = '{87.2253352734, -71.4507268762, -76.4236341226, 28.7819654885, 83.650076119, 61.8395212632, 62.1094886394, -27.9292168869};
test_label[2295] = '{87.2253352734};
test_output[2295] = '{0.0276231109876};
############ END DEBUG ############*/
test_input[18368:18375] = '{32'hc150d68a, 32'h426afb17, 32'hc164e5d2, 32'hc252baa4, 32'hc293027a, 32'h41b6cde5, 32'h4226917a, 32'hc1df5ff3};
test_label[2296] = '{32'hc252baa4};
test_output[2296] = '{32'h42dedade};
/*############ DEBUG ############
test_input[18368:18375] = '{-13.0523775701, 58.7452049289, -14.3061082014, -52.6822662751, -73.5048402552, 22.8505352111, 41.6420681161, -27.9218502081};
test_label[2296] = '{-52.6822662751};
test_output[2296] = '{111.427471241};
############ END DEBUG ############*/
test_input[18376:18383] = '{32'hc20cd337, 32'h414e8a70, 32'hc25ab2c0, 32'hc21dfaf2, 32'hc2b33ac4, 32'hc2a7de42, 32'hc2803165, 32'hc23ecf10};
test_label[2297] = '{32'hc2b33ac4};
test_output[2297] = '{32'h42cd0c12};
/*############ DEBUG ############
test_input[18376:18383] = '{-35.206262698, 12.9087986749, -54.6745594838, -39.495065135, -89.6147773967, -83.9341000581, -64.096472246, -47.7022088148};
test_label[2297] = '{-89.6147773967};
test_output[2297] = '{102.523576072};
############ END DEBUG ############*/
test_input[18384:18391] = '{32'h42553455, 32'hc2a12685, 32'hc0a6be3f, 32'h42c011ca, 32'h42684cd8, 32'hc237945a, 32'h4205412c, 32'h42ada677};
test_label[2298] = '{32'h4205412c};
test_output[2298] = '{32'h427ae282};
/*############ DEBUG ############
test_input[18384:18391] = '{53.301104709, -80.5752329133, -5.21072324645, 96.0347413015, 58.0750442591, -45.8948738589, 33.3136440912, 86.8251292242};
test_label[2298] = '{33.3136440912};
test_output[2298] = '{62.7211972782};
############ END DEBUG ############*/
test_input[18392:18399] = '{32'hc2becca4, 32'h41edf862, 32'h4121b1a4, 32'h41415e01, 32'h42bf5c5a, 32'hc214ba58, 32'h41c917b2, 32'hc250d07f};
test_label[2299] = '{32'hc214ba58};
test_output[2299] = '{32'h4304dcc3};
/*############ DEBUG ############
test_input[18392:18399] = '{-95.3996849985, 29.7462813933, 10.1058694166, 12.0854505855, 95.6803735091, -37.1819780045, 25.1365693032, -52.203609181};
test_label[2299] = '{-37.1819780045};
test_output[2299] = '{132.862351514};
############ END DEBUG ############*/
test_input[18400:18407] = '{32'h4235ed7b, 32'h429cbba3, 32'hc1d76cec, 32'hc0291b66, 32'hc2b48b13, 32'h4152c7bb, 32'h427a54b5, 32'h42a89f70};
test_label[2300] = '{32'h4152c7bb};
test_output[2300] = '{32'h428e47cf};
/*############ DEBUG ############
test_input[18400:18407] = '{45.481916134, 78.3664798953, -26.9281835947, -2.64229734652, -90.2716324646, 13.1737625908, 62.5827220075, 84.3113992956};
test_label[2300] = '{13.1737625908};
test_output[2300] = '{71.1402523947};
############ END DEBUG ############*/
test_input[18408:18415] = '{32'hc210d71a, 32'hc24b7ba3, 32'hc2448a2a, 32'h427942c5, 32'hc263db6e, 32'h428dcdc0, 32'h4193c044, 32'h42959eab};
test_label[2301] = '{32'h428dcdc0};
test_output[2301] = '{32'h407b631b};
/*############ DEBUG ############
test_input[18408:18415] = '{-36.2100614194, -50.8707375768, -49.1349258906, 62.3152048955, -56.964286563, 70.9018556976, 18.4688805047, 74.809894978};
test_label[2301] = '{70.9018556976};
test_output[2301] = '{3.92792384543};
############ END DEBUG ############*/
test_input[18416:18423] = '{32'hc2c49171, 32'hc2b391f7, 32'h414c97b1, 32'hc27ffa89, 32'h41ce01fc, 32'hc1d8547c, 32'h4166edfa, 32'hc2851419};
test_label[2302] = '{32'hc2851419};
test_output[2302] = '{32'h42b8949a};
/*############ DEBUG ############
test_input[18416:18423] = '{-98.2840639231, -89.7850867499, 12.7870344766, -63.9946626656, 25.7509681412, -27.0412527029, 14.4330996255, -66.5392512617};
test_label[2302] = '{-66.5392512617};
test_output[2302] = '{92.2902338999};
############ END DEBUG ############*/
test_input[18424:18431] = '{32'hc2a556c7, 32'h42a69e93, 32'h4245c87a, 32'hc2c66a5f, 32'hc2aef6d0, 32'h420f511b, 32'hc1f8c01b, 32'hc229b92b};
test_label[2303] = '{32'hc2a556c7};
test_output[2303] = '{32'h4325faad};
/*############ DEBUG ############
test_input[18424:18431] = '{-82.6694838854, 83.3097187818, 49.4457788214, -99.2077588666, -87.4820588447, 35.8292043101, -31.0938017726, -42.4308286351};
test_label[2303] = '{-82.6694838854};
test_output[2303] = '{165.979202667};
############ END DEBUG ############*/
test_input[18432:18439] = '{32'h42a8a937, 32'h42b4c8be, 32'h42bce367, 32'h42802293, 32'h425373c0, 32'hc1c5d955, 32'h42a1f1ef, 32'hc2b19d78};
test_label[2304] = '{32'h42bce367};
test_output[2304] = '{32'h3c8d8ae9};
/*############ DEBUG ############
test_input[18432:18439] = '{84.3304963298, 90.3920750835, 94.4441450166, 64.0675289881, 52.8630379644, -24.7311198848, 80.9725279348, -88.8075567995};
test_label[2304] = '{94.4441450166};
test_output[2304] = '{0.0172781512288};
############ END DEBUG ############*/
test_input[18440:18447] = '{32'h41fbed08, 32'hc210b396, 32'h4283415e, 32'h4217c06a, 32'h4255a0de, 32'h42611c54, 32'h42bb929c, 32'hc2b49baf};
test_label[2305] = '{32'h42611c54};
test_output[2305] = '{32'h421608e5};
/*############ DEBUG ############
test_input[18440:18447] = '{31.4907387371, -36.1753762707, 65.6276733435, 37.9379034462, 53.407095096, 56.2776631781, 93.7863482766, -90.3040701022};
test_label[2305] = '{56.2776631781};
test_output[2305] = '{37.5086850985};
############ END DEBUG ############*/
test_input[18448:18455] = '{32'hbff140ac, 32'h41d73f06, 32'hc23b64ec, 32'hc272ac2d, 32'h429e9c1d, 32'hc20001db, 32'h4215e311, 32'hc142967d};
test_label[2306] = '{32'h4215e311};
test_output[2306] = '{32'h42275529};
/*############ DEBUG ############
test_input[18448:18455] = '{-1.88478615693, 26.9057727308, -46.8485558602, -60.6681398684, 79.3049103226, -32.0018104201, 37.4717450044, -12.1617404054};
test_label[2306] = '{37.4717450044};
test_output[2306] = '{41.8331653181};
############ END DEBUG ############*/
test_input[18456:18463] = '{32'hc2c73b5b, 32'h3ff89f64, 32'hc25a3168, 32'hc223e8b3, 32'hc289818b, 32'hc24ac6f3, 32'hc1ee3098, 32'hc299a453};
test_label[2307] = '{32'hc1ee3098};
test_output[2307] = '{32'h41fdba8e};
/*############ DEBUG ############
test_input[18456:18463] = '{-99.6159321968, 1.94236416174, -54.5482500761, -40.9772466268, -68.7530149756, -50.6942851516, -29.7737268467, -76.8209428145};
test_label[2307] = '{-29.7737268467};
test_output[2307] = '{31.7160910084};
############ END DEBUG ############*/
test_input[18464:18471] = '{32'h4231424e, 32'h42aad7be, 32'h42994b63, 32'h41f1d17d, 32'h4154bf94, 32'hc16d0e85, 32'hc1d39e17, 32'h421b7240};
test_label[2308] = '{32'h4154bf94};
test_output[2308] = '{32'h42903fe0};
/*############ DEBUG ############
test_input[18464:18471] = '{44.3147520301, 85.4213734963, 76.6472386971, 30.2272883209, 13.2967723096, -14.8160447389, -26.452191376, 38.861574057};
test_label[2308] = '{13.2967723096};
test_output[2308] = '{72.1247558574};
############ END DEBUG ############*/
test_input[18472:18479] = '{32'hc2aedaf0, 32'hc2873e7a, 32'h4222542d, 32'h429a7823, 32'h420391c2, 32'hc18bdef8, 32'h419d0e92, 32'hc1cf4900};
test_label[2309] = '{32'hc1cf4900};
test_output[2309] = '{32'h42ce4a63};
/*############ DEBUG ############
test_input[18472:18479] = '{-87.4276134432, -67.6220247478, 40.5822027086, 77.2346401999, 32.8923433308, -17.483870594, 19.632114561, -25.9106449805};
test_label[2309] = '{-25.9106449805};
test_output[2309] = '{103.14528518};
############ END DEBUG ############*/
test_input[18480:18487] = '{32'hc280ad69, 32'hc233b1fc, 32'hc1fb16b3, 32'h41c2825b, 32'hc221969f, 32'h4212d45f, 32'hc251b939, 32'hc29adda5};
test_label[2310] = '{32'hc221969f};
test_output[2310] = '{32'h429a3580};
/*############ DEBUG ############
test_input[18480:18487] = '{-64.338690763, -44.9238137093, -31.386083925, 24.3136503439, -40.3970927329, 36.7073948274, -52.4308824705, -77.4328971328};
test_label[2310] = '{-40.3970927329};
test_output[2310] = '{77.1044917047};
############ END DEBUG ############*/
test_input[18488:18495] = '{32'hc2bda38d, 32'h428eefe5, 32'h429639f6, 32'h42b39412, 32'hc2a376a9, 32'h4221f72d, 32'hc27b85a1, 32'h41f09dbd};
test_label[2311] = '{32'h429639f6};
test_output[2311] = '{32'h416ad0dd};
/*############ DEBUG ############
test_input[18488:18495] = '{-94.819432271, 71.4685412671, 75.1132075236, 89.7891988481, -81.7317577928, 40.4913813664, -62.8804983918, 30.0770201371};
test_label[2311] = '{75.1132075236};
test_output[2311] = '{14.6759917585};
############ END DEBUG ############*/
test_input[18496:18503] = '{32'h429d1e42, 32'hc1edc100, 32'hc2afa12e, 32'hc282563f, 32'h42b42c1d, 32'hc284840a, 32'h427dd1bc, 32'hc211a5b9};
test_label[2312] = '{32'h429d1e42};
test_output[2312] = '{32'h41386ee9};
/*############ DEBUG ############
test_input[18496:18503] = '{78.5590936297, -29.7192381636, -87.814802129, -65.1684513451, 90.0861610187, -66.25788888, 63.4548186545, -36.4118381245};
test_label[2312] = '{78.5590936297};
test_output[2312] = '{11.5270772485};
############ END DEBUG ############*/
test_input[18504:18511] = '{32'h422fe01e, 32'h41bb7a17, 32'hc2a1b55a, 32'h40172820, 32'hc2bd574c, 32'hc215694f, 32'h42a78f2c, 32'hc17bc4a6};
test_label[2313] = '{32'hc2bd574c};
test_output[2313] = '{32'h4332733c};
/*############ DEBUG ############
test_input[18504:18511] = '{43.9688650275, 23.4346139145, -80.8541984753, 2.36182407635, -94.6705013362, -37.3528390581, 83.7796302365, -15.7355098274};
test_label[2313] = '{-94.6705013362};
test_output[2313] = '{178.450131573};
############ END DEBUG ############*/
test_input[18512:18519] = '{32'h42a56d01, 32'h421ab56a, 32'h42c0fd61, 32'h42a88558, 32'h411a0a3b, 32'h41479eae, 32'hc0c75abe, 32'h42611deb};
test_label[2314] = '{32'h42c0fd61};
test_output[2314] = '{32'h36c5c6ca};
/*############ DEBUG ############
test_input[18512:18519] = '{82.7128999422, 38.677162925, 96.4948827491, 84.2604355153, 9.62749747347, 12.4762403062, -6.22982672819, 56.2792165177};
test_label[2314] = '{96.4948827491};
test_output[2314] = '{5.89419971852e-06};
############ END DEBUG ############*/
test_input[18520:18527] = '{32'hc2c6d20e, 32'hc1ed66f3, 32'hc22cfe01, 32'hc17f9f9e, 32'h42b6621e, 32'hc290efe3, 32'h42ab30e1, 32'hc1864ebc};
test_label[2315] = '{32'hc17f9f9e};
test_output[2315] = '{32'h42d657f7};
/*############ DEBUG ############
test_input[18520:18527] = '{-99.4102593799, -29.6752676274, -43.2480524875, -15.9764692776, 91.1916348941, -72.4685298682, 85.5954655841, -16.7884435828};
test_label[2315] = '{-15.9764692776};
test_output[2315] = '{107.171809355};
############ END DEBUG ############*/
test_input[18528:18535] = '{32'h42a8ad74, 32'hc1d51604, 32'hc0f79de1, 32'h418ab287, 32'hc1a1daf2, 32'h41d3a72e, 32'hc29bc961, 32'hc29451eb};
test_label[2316] = '{32'h41d3a72e};
test_output[2316] = '{32'h42678751};
/*############ DEBUG ############
test_input[18528:18535] = '{84.3387738477, -26.6357496157, -7.73802242183, 17.3371719505, -20.2319074495, 26.4566299315, -77.893318665, -74.1599967293};
test_label[2316] = '{26.4566299315};
test_output[2316] = '{57.8821439162};
############ END DEBUG ############*/
test_input[18536:18543] = '{32'h41cb93af, 32'h42117b5b, 32'hc2832b20, 32'h428cd3e5, 32'hc2a40024, 32'hc25b7287, 32'hc238dae5, 32'h42606c0c};
test_label[2317] = '{32'h42117b5b};
test_output[2317] = '{32'h42082c6f};
/*############ DEBUG ############
test_input[18536:18543] = '{25.4471119086, 36.370465593, -65.5842307717, 70.4138562555, -82.0002756049, -54.8618448369, -46.2137658268, 56.1055154649};
test_label[2317] = '{36.370465593};
test_output[2317] = '{34.0433912734};
############ END DEBUG ############*/
test_input[18544:18551] = '{32'h42afa2ab, 32'h3e9199bf, 32'hc279709b, 32'hc11b6ec1, 32'h42c4c888, 32'h41f577d3, 32'h41b189a3, 32'h3fc70ef2};
test_label[2318] = '{32'h41b189a3};
test_output[2318] = '{32'h42986623};
/*############ DEBUG ############
test_input[18544:18551] = '{87.8177138253, 0.284376112009, -62.3599671526, -9.71453966372, 98.3916655107, 30.6835075304, 22.1922055752, 1.55514364558};
test_label[2318] = '{22.1922055752};
test_output[2318] = '{76.1994855088};
############ END DEBUG ############*/
test_input[18552:18559] = '{32'hc1843d53, 32'h40c81b2c, 32'hc17c3dac, 32'hc259e58b, 32'h420c278c, 32'hc0910428, 32'hc232e317, 32'hc2058366};
test_label[2319] = '{32'hc17c3dac};
test_output[2319] = '{32'h424b36f7};
/*############ DEBUG ############
test_input[18552:18559] = '{-16.5299425885, 6.25331667987, -15.7650570108, -54.4741621599, 35.0386210373, -4.53175755598, -44.721766957, -33.3783179764};
test_label[2319] = '{-15.7650570108};
test_output[2319] = '{50.8036780481};
############ END DEBUG ############*/
test_input[18560:18567] = '{32'hc127dd25, 32'h42b0d387, 32'hc28e27f4, 32'h421e8fc5, 32'h4288a993, 32'hc2299809, 32'hc28fa872, 32'h40746dc8};
test_label[2320] = '{32'hc2299809};
test_output[2320] = '{32'h4302cfc6};
/*############ DEBUG ############
test_input[18560:18567] = '{-10.4914902713, 88.4131412572, -71.0780372245, 39.6403987815, 68.3311965779, -42.3984708441, -71.828993668, 3.81920057194};
test_label[2320] = '{-42.3984708441};
test_output[2320] = '{130.811612103};
############ END DEBUG ############*/
test_input[18568:18575] = '{32'h40e77d9d, 32'h3ffe75bf, 32'hc11da0f0, 32'hc296859d, 32'h40ba79e7, 32'hc1b80a17, 32'h415bbb0c, 32'h41c31ecf};
test_label[2321] = '{32'h3ffe75bf};
test_output[2321] = '{32'h41b3377f};
/*############ DEBUG ############
test_input[18568:18575] = '{7.23408372329, 1.98796830042, -9.85179137215, -75.2609631297, 5.82738057899, -23.0049258447, 13.7331660275, 24.3900425353};
test_label[2321] = '{1.98796830042};
test_output[2321] = '{22.4020978173};
############ END DEBUG ############*/
test_input[18576:18583] = '{32'h415a388d, 32'hbf3a06fa, 32'h42177354, 32'h41b345a4, 32'h428dd3db, 32'hc2a4aca7, 32'hc0f535d8, 32'hc2339274};
test_label[2322] = '{32'h41b345a4};
test_output[2322] = '{32'h424204e4};
/*############ DEBUG ############
test_input[18576:18583] = '{13.6388060812, -0.726668970798, 37.8626245767, 22.409003417, 70.9137780941, -82.337215273, -7.66282262098, -44.8930211369};
test_label[2322] = '{22.409003417};
test_output[2322] = '{48.5047746771};
############ END DEBUG ############*/
test_input[18584:18591] = '{32'hc285584b, 32'h429714cc, 32'h41d80dc6, 32'h4133a4ec, 32'h41d71b4b, 32'h41e5a317, 32'hc226fa33, 32'hc1b9b556};
test_label[2323] = '{32'hc226fa33};
test_output[2323] = '{32'h42ea91e6};
/*############ DEBUG ############
test_input[18584:18591] = '{-66.6724478436, 75.5406199303, 27.0067262287, 11.2277640423, 26.888325957, 28.7046336482, -41.744336444, -23.2135436613};
test_label[2323] = '{-41.744336444};
test_output[2323] = '{117.284956374};
############ END DEBUG ############*/
test_input[18592:18599] = '{32'h423a9a4d, 32'hc18f6e5d, 32'hc28802b2, 32'h42a81db9, 32'hc20b6569, 32'h415d017d, 32'hc187b32a, 32'hc2c33e61};
test_label[2324] = '{32'h415d017d};
test_output[2324] = '{32'h428c7d8a};
/*############ DEBUG ############
test_input[18592:18599] = '{46.6506827645, -17.9288888364, -68.0052662528, 84.0580549405, -34.8490337536, 13.8128636337, -16.9624834039, -97.6218333793};
test_label[2324] = '{13.8128636337};
test_output[2324] = '{70.2451913068};
############ END DEBUG ############*/
test_input[18600:18607] = '{32'h42c01026, 32'h422d2479, 32'h42a2b03f, 32'h40442c7c, 32'hc2918d9c, 32'h42712def, 32'h40845fce, 32'hc1992b79};
test_label[2325] = '{32'h42a2b03f};
test_output[2325] = '{32'h416aff39};
/*############ DEBUG ############
test_input[18600:18607] = '{96.031543373, 43.2856175068, 81.3442334118, 3.06521513897, -72.7765816335, 60.2948567672, 4.13669505804, -19.1462272371};
test_label[2325] = '{81.3442334118};
test_output[2325] = '{14.6873103794};
############ END DEBUG ############*/
test_input[18608:18615] = '{32'h402fd0f0, 32'hc2316221, 32'h41afface, 32'hc10f7227, 32'h42a9cb35, 32'hc258ca8c, 32'hc214311c, 32'h41e7e706};
test_label[2326] = '{32'hc258ca8c};
test_output[2326] = '{32'h430b183e};
/*############ DEBUG ############
test_input[18608:18615] = '{2.74712750252, -44.3458288565, 21.9974625982, -8.96536885318, 84.8968902304, -54.1978013517, -37.047958782, 28.9878034891};
test_label[2326] = '{-54.1978013517};
test_output[2326] = '{139.094691582};
############ END DEBUG ############*/
test_input[18616:18623] = '{32'h4279d1f7, 32'hc293611a, 32'h42107e94, 32'hc225118f, 32'hc1e44530, 32'hc1a18805, 32'hc25f9b78, 32'h422e27a2};
test_label[2327] = '{32'hc293611a};
test_output[2327] = '{32'h4308250b};
/*############ DEBUG ############
test_input[18616:18623] = '{62.4550456812, -73.6896522305, 36.1236100974, -41.2671475111, -28.5337820676, -20.1914154913, -55.9018231506, 43.5387046967};
test_label[2327] = '{-73.6896522305};
test_output[2327] = '{136.144697918};
############ END DEBUG ############*/
test_input[18624:18631] = '{32'hc2126086, 32'hc1a53976, 32'h41b7f14e, 32'hc244b280, 32'h42879701, 32'hc2c66255, 32'h4239b85a, 32'hc1babe82};
test_label[2328] = '{32'h4239b85a};
test_output[2328] = '{32'h41aaeb50};
/*############ DEBUG ############
test_input[18624:18631] = '{-36.5942603119, -20.65305704, 22.9928239177, -49.1743148586, 67.7949309389, -99.1920553299, 46.430031709, -23.3430219842};
test_label[2328] = '{46.430031709};
test_output[2328] = '{21.3648992304};
############ END DEBUG ############*/
test_input[18632:18639] = '{32'hc20d25a7, 32'h42682ad4, 32'hc2053a2d, 32'hc29a4c8d, 32'h422ccf39, 32'h42ac82c6, 32'hc290e5e4, 32'h42954277};
test_label[2329] = '{32'hc29a4c8d};
test_output[2329] = '{32'h432367aa};
/*############ DEBUG ############
test_input[18632:18639] = '{-35.2867694753, 58.0418237456, -33.306811225, -77.1495134459, 43.2023649814, 86.2554181033, -72.4490089324, 74.6298124906};
test_label[2329] = '{-77.1495134459};
test_output[2329] = '{163.404940484};
############ END DEBUG ############*/
test_input[18640:18647] = '{32'h42a27608, 32'h42ab0ce0, 32'hc2a712ff, 32'h41cc7b86, 32'hc1924565, 32'h4196e43a, 32'hc2ba32d4, 32'h4147c140};
test_label[2330] = '{32'hc1924565};
test_output[2330] = '{32'h42cfa529};
/*############ DEBUG ############
test_input[18640:18647] = '{81.2305272461, 85.5251453547, -83.5371034461, 25.5603137752, -18.2838833686, 18.8614386505, -93.0992718137, 12.4846801634};
test_label[2330] = '{-18.2838833686};
test_output[2330] = '{103.822578292};
############ END DEBUG ############*/
test_input[18648:18655] = '{32'h423714ab, 32'hc2c6654e, 32'hc27b4cb9, 32'hc2b35bd0, 32'hc115b6b4, 32'hc28cbf06, 32'h40144816, 32'hc2b13f3d};
test_label[2331] = '{32'hc2c6654e};
test_output[2331] = '{32'h4310f7d2};
/*############ DEBUG ############
test_input[18648:18655] = '{45.7701836019, -99.1978586403, -62.8249238638, -89.6793195416, -9.35710544055, -70.3730903873, 2.31689970101, -88.6235131312};
test_label[2331] = '{-99.1978586403};
test_output[2331] = '{144.968042242};
############ END DEBUG ############*/
test_input[18656:18663] = '{32'h41a25a5a, 32'h41490fe9, 32'h4220c783, 32'h426e5923, 32'h42672672, 32'h4222a3c8, 32'hc217160e, 32'h42b8c175};
test_label[2332] = '{32'hc217160e};
test_output[2332] = '{32'h4302263e};
/*############ DEBUG ############
test_input[18656:18663] = '{20.2941175843, 12.5663844294, 40.1948345019, 59.5870458819, 57.7875456959, 40.6599417818, -37.7715364322, 92.3778426652};
test_label[2332] = '{-37.7715364322};
test_output[2332] = '{130.149379097};
############ END DEBUG ############*/
test_input[18664:18671] = '{32'hc1c675c1, 32'h422c3f11, 32'hc1d27a22, 32'h42b739cd, 32'h42c53ee5, 32'hc1806587, 32'h4191419d, 32'hc19741cd};
test_label[2333] = '{32'h422c3f11};
test_output[2333] = '{32'h425e3fa5};
/*############ DEBUG ############
test_input[18664:18671] = '{-24.807497721, 43.0615894708, -26.309635241, 91.6128921932, 98.6228402069, -16.0495742176, 18.1570380721, -18.9071290678};
test_label[2333] = '{43.0615894708};
test_output[2333] = '{55.5621531844};
############ END DEBUG ############*/
test_input[18672:18679] = '{32'hc2a6e85b, 32'h428fae9d, 32'hbd97fc23, 32'hc27128a4, 32'hc2a69d40, 32'h41ffb66f, 32'hc2642029, 32'h428e6d2f};
test_label[2334] = '{32'hc2642029};
test_output[2334] = '{32'h43014cd8};
/*############ DEBUG ############
test_input[18672:18679] = '{-83.4538170382, 71.8410401435, -0.0742113842968, -60.2896881263, -83.3071304379, 31.9640784273, -57.0314080296, 71.2132455296};
test_label[2334] = '{-57.0314080296};
test_output[2334] = '{129.300175409};
############ END DEBUG ############*/
test_input[18680:18687] = '{32'hc1c4cd12, 32'h41f96df1, 32'hc2749137, 32'h42b29f12, 32'h41ab869a, 32'hc250052d, 32'h42972eb8, 32'h3ffe5b5e};
test_label[2335] = '{32'h3ffe5b5e};
test_output[2335] = '{32'h42aea5a5};
/*############ DEBUG ############
test_input[18680:18687] = '{-24.6001311846, 31.178683186, -61.1418119908, 89.3106866827, 21.4407234168, -52.0050557925, 75.5912452601, 1.98716333534};
test_label[2335] = '{1.98716333534};
test_output[2335] = '{87.3235244482};
############ END DEBUG ############*/
test_input[18688:18695] = '{32'h41e45c83, 32'h415e5ba3, 32'hc2bc6697, 32'hc18c1f75, 32'h42666c13, 32'hc242d97a, 32'hc1326731, 32'h4219df76};
test_label[2336] = '{32'hc242d97a};
test_output[2336] = '{32'h42d4a2c7};
/*############ DEBUG ############
test_input[18688:18695] = '{28.5451712792, 13.8973725577, -94.2003671566, -17.5153606055, 57.6055430826, -48.712380806, -11.1501935474, 38.468222458};
test_label[2336] = '{-48.712380806};
test_output[2336] = '{106.317923893};
############ END DEBUG ############*/
test_input[18696:18703] = '{32'h419e0755, 32'hc10bf3b0, 32'h428d78e5, 32'h4076c5e9, 32'h426df537, 32'h41d64482, 32'h428aded0, 32'h41fb11c8};
test_label[2337] = '{32'h419e0755};
test_output[2337] = '{32'h424ce4b9};
/*############ DEBUG ############
test_input[18696:18703] = '{19.7535795959, -8.74699429756, 70.7361249326, 3.85582940157, 59.4894691594, 26.7834517366, 69.4351806192, 31.3836828866};
test_label[2337] = '{19.7535795959};
test_output[2337] = '{51.2233618845};
############ END DEBUG ############*/
test_input[18704:18711] = '{32'hc2ba2d21, 32'h424c2611, 32'h42098f4b, 32'hc29071a6, 32'h4286bea8, 32'h3f88cb6a, 32'h42a73795, 32'h4280026b};
test_label[2338] = '{32'h4280026b};
test_output[2338] = '{32'h419cd4a9};
/*############ DEBUG ############
test_input[18704:18711] = '{-93.0881459524, 51.0371727265, 34.3899345861, -72.2219706922, 67.3723732674, 1.06870774583, 83.6085609309, 64.0047238682};
test_label[2338] = '{64.0047238682};
test_output[2338] = '{19.6038371546};
############ END DEBUG ############*/
test_input[18712:18719] = '{32'h42829077, 32'h3fa13db1, 32'h41c04479, 32'hc1f67208, 32'hc2074902, 32'hc23eddbf, 32'h4221858b, 32'hc297ba64};
test_label[2339] = '{32'hc2074902};
test_output[2339] = '{32'h42c634f8};
/*############ DEBUG ############
test_input[18712:18719] = '{65.2821569402, 1.25969517221, 24.0334333162, -30.8056790533, -33.82129806, -47.7165497086, 40.3804131712, -75.8640428152};
test_label[2339] = '{-33.82129806};
test_output[2339] = '{99.1034550003};
############ END DEBUG ############*/
test_input[18720:18727] = '{32'hc23f2ec9, 32'hc26936ef, 32'h4288a31a, 32'h42239f65, 32'h429196d2, 32'hc28dca18, 32'hc2731412, 32'h41944598};
test_label[2340] = '{32'hc26936ef};
test_output[2340] = '{32'h43031c0a};
/*############ DEBUG ############
test_input[18720:18727] = '{-47.7956869977, -58.3036450324, 68.3185597157, 40.9056601121, 72.7945740333, -70.8947109976, -60.769599163, 18.5339810759};
test_label[2340] = '{-58.3036450324};
test_output[2340] = '{131.10953349};
############ END DEBUG ############*/
test_input[18728:18735] = '{32'hc21a752f, 32'h429d94e9, 32'h417fa1db, 32'h420854cd, 32'h423da670, 32'h41d9a780, 32'h4292150a, 32'h41fbeb83};
test_label[2341] = '{32'h4292150a};
test_output[2341] = '{32'h40b817f9};
/*############ DEBUG ############
test_input[18728:18735] = '{-38.6144352339, 78.7908381468, 15.9770157305, 34.0828125656, 47.412536461, 27.2067869866, 73.0410901593, 31.4899961003};
test_label[2341] = '{73.0410901593};
test_output[2341] = '{5.7529265137};
############ END DEBUG ############*/
test_input[18736:18743] = '{32'h4134a482, 32'hc2868d81, 32'h41986f85, 32'hc1a47dea, 32'hc2c32372, 32'h427c8468, 32'h42a10f41, 32'hc0ce17ef};
test_label[2342] = '{32'hc0ce17ef};
test_output[2342] = '{32'h42adf0c0};
/*############ DEBUG ############
test_input[18736:18743] = '{11.2901627099, -67.2763737589, 19.0544521899, -20.5614811999, -97.5692296915, 63.1293013606, 80.5297943826, -6.44042134802};
test_label[2342] = '{-6.44042134802};
test_output[2342] = '{86.9702157584};
############ END DEBUG ############*/
test_input[18744:18751] = '{32'hc01776a4, 32'hc2beb53f, 32'h40c8f93d, 32'hc1e46a10, 32'h4255e4c9, 32'h41bdf41b, 32'hc29b83da, 32'h42521999};
test_label[2343] = '{32'hc01776a4};
test_output[2343] = '{32'h4260ab74};
/*############ DEBUG ############
test_input[18744:18751] = '{-2.36661627999, -95.3539940278, 6.28042445518, -28.5517879476, 53.4734233762, 23.7441925619, -77.7575212614, 52.5249994695};
test_label[2343] = '{-2.36661627999};
test_output[2343] = '{56.1674358614};
############ END DEBUG ############*/
test_input[18752:18759] = '{32'h429bb010, 32'hc2a6d77b, 32'hc2aa6eed, 32'hc29c6252, 32'h42b423cf, 32'h42a1c4e2, 32'hc117b54a, 32'h42287bf4};
test_label[2344] = '{32'hc2aa6eed};
test_output[2344] = '{32'h432f4965};
/*############ DEBUG ############
test_input[18752:18759] = '{77.8438741722, -83.4208567449, -85.2166555998, -78.1920300927, 90.0699407983, 80.8845345308, -9.48176043923, 42.1210473338};
test_label[2344] = '{-85.2166555998};
test_output[2344] = '{175.286703818};
############ END DEBUG ############*/
test_input[18760:18767] = '{32'h4290fab5, 32'hc1a3b5d7, 32'hc0b92197, 32'hc29c31bc, 32'h429de074, 32'hc2636ba2, 32'hc27e0c2e, 32'hc29f5375};
test_label[2345] = '{32'h4290fab5};
test_output[2345] = '{32'h40ce68e7};
/*############ DEBUG ############
test_input[18760:18767] = '{72.4896624653, -20.4637892139, -5.78535025626, -78.0971379567, 78.9383866551, -56.8551083543, -63.5118950865, -79.663003286};
test_label[2345] = '{72.4896624653};
test_output[2345] = '{6.45030547879};
############ END DEBUG ############*/
test_input[18768:18775] = '{32'h41ce1997, 32'h421d74b9, 32'hc04def3a, 32'h4216b5f1, 32'hc2285d3e, 32'hc28b6b2b, 32'h422dfe51, 32'h4197723a};
test_label[2346] = '{32'hc04def3a};
test_output[2346] = '{32'h423af085};
/*############ DEBUG ############
test_input[18768:18775] = '{25.7624942802, 39.3639880974, -3.2177262533, 37.677677667, -42.0910581783, -69.7093104593, 43.4983547818, 18.9307750831};
test_label[2346] = '{-3.2177262533};
test_output[2346] = '{46.7348816108};
############ END DEBUG ############*/
test_input[18776:18783] = '{32'hc10c73ff, 32'h41f1e1e0, 32'hc10ccadb, 32'hc2557f91, 32'h421ef38a, 32'hc205a013, 32'hc1e0804c, 32'h42ac2633};
test_label[2347] = '{32'hc10c73ff};
test_output[2347] = '{32'h42bdb4b3};
/*############ DEBUG ############
test_input[18776:18783] = '{-8.77831895684, 30.2352899226, -8.79952522582, -53.3745766937, 39.737830686, -33.4063211952, -28.0626453971, 86.0746078829};
test_label[2347] = '{-8.77831895684};
test_output[2347] = '{94.8529268398};
############ END DEBUG ############*/
test_input[18784:18791] = '{32'hc1c1bd45, 32'hc239f83f, 32'hc2a629d3, 32'h42baf2da, 32'hc238d47d, 32'h42340240, 32'h429927b9, 32'hc26dbbc3};
test_label[2348] = '{32'hc26dbbc3};
test_output[2348] = '{32'h4318e85e};
/*############ DEBUG ############
test_input[18784:18791] = '{-24.217417282, -46.4924287013, -83.0816911841, 93.4743221698, -46.2075064067, 45.00219646, 76.5775799975, -59.4333614247};
test_label[2348] = '{-59.4333614247};
test_output[2348] = '{152.90768364};
############ END DEBUG ############*/
test_input[18792:18799] = '{32'h429f3d13, 32'h4258bcf1, 32'hc1dd0681, 32'hc1ace34e, 32'h42aece4c, 32'hc276b057, 32'h42344a7e, 32'h412799eb};
test_label[2349] = '{32'hc1dd0681};
test_output[2349] = '{32'h42e61023};
/*############ DEBUG ############
test_input[18792:18799] = '{79.6192826359, 54.184511575, -27.6281765738, -21.6109886426, 87.4029215484, -61.6722080158, 45.07274668, 10.4750775744};
test_label[2349] = '{-27.6281765738};
test_output[2349] = '{115.031514529};
############ END DEBUG ############*/
test_input[18800:18807] = '{32'h42a491ea, 32'hc194d2a3, 32'h42a507df, 32'h424487b7, 32'hc1c4933d, 32'hc28d994e, 32'h4290c617, 32'hc298f83d};
test_label[2350] = '{32'h42a507df};
test_output[2350] = '{32'h3f15a7f2};
/*############ DEBUG ############
test_input[18800:18807] = '{82.2849848255, -18.6028507372, 82.5153768182, 49.1325343706, -24.5718935696, -70.7994238327, 72.3868941212, -76.4848372888};
test_label[2350] = '{82.5153768182};
test_output[2350] = '{0.584593872344};
############ END DEBUG ############*/
test_input[18808:18815] = '{32'h42112ce0, 32'hc2320972, 32'hc1d1d453, 32'hc256f501, 32'hc2b3f9ab, 32'h41f875d9, 32'h418949f9, 32'hc29a9458};
test_label[2351] = '{32'h41f875d9};
test_output[2351] = '{32'h40a7bb13};
/*############ DEBUG ############
test_input[18808:18815] = '{36.2938225604, -44.5092247774, -26.2286730469, -53.7392608463, -89.9876353904, 31.0575423078, 17.1611203585, -77.2897305553};
test_label[2351] = '{31.0575423078};
test_output[2351] = '{5.24158616539};
############ END DEBUG ############*/
test_input[18816:18823] = '{32'h42b1ecbd, 32'hc2baf764, 32'hc13302ca, 32'h429d0642, 32'hc1c46252, 32'h4270967b, 32'hc2b82334, 32'h41fb008c};
test_label[2352] = '{32'hc2b82334};
test_output[2352] = '{32'h433507fa};
/*############ DEBUG ############
test_input[18816:18823] = '{88.9623761715, -93.4831838297, -11.1881808715, 78.5122210059, -24.5480087243, 60.1469528453, -92.0687525, 31.3752678191};
test_label[2352] = '{-92.0687525};
test_output[2352] = '{181.031157615};
############ END DEBUG ############*/
test_input[18824:18831] = '{32'h416b7643, 32'hc25f365f, 32'h4297cd2b, 32'hc06618b2, 32'hc2a2eb30, 32'hc24ec2a5, 32'h420fca21, 32'hc28a19f8};
test_label[2353] = '{32'hc28a19f8};
test_output[2353] = '{32'h4310f391};
/*############ DEBUG ############
test_input[18824:18831] = '{14.7163727546, -55.8030966063, 75.9007180161, -3.59525729415, -81.459349116, -51.6900829825, 35.947390386, -69.0507198972};
test_label[2353] = '{-69.0507198972};
test_output[2353] = '{144.951437913};
############ END DEBUG ############*/
test_input[18832:18839] = '{32'h42960cdc, 32'hc2a2cf6c, 32'hc200cb92, 32'h428c567f, 32'h42a35be4, 32'hc274e32f, 32'h42aa6699, 32'hc1e24a38};
test_label[2354] = '{32'hc274e32f};
test_output[2354] = '{32'h43127391};
/*############ DEBUG ############
test_input[18832:18839] = '{75.0251179408, -81.4051226962, -32.1987986514, 70.1689375236, 81.6794728379, -61.2218594569, 85.2003847852, -28.2862387258};
test_label[2354] = '{-61.2218594569};
test_output[2354] = '{146.451425159};
############ END DEBUG ############*/
test_input[18840:18847] = '{32'hc2029ceb, 32'hc27b9611, 32'h42a94e06, 32'hc001009e, 32'hc294040a, 32'hc14905a6, 32'h42812fe0, 32'hbf0015cd};
test_label[2355] = '{32'h42812fe0};
test_output[2355] = '{32'h41a07897};
/*############ DEBUG ############
test_input[18840:18847] = '{-32.6532392837, -62.8965478098, 84.6523880959, -2.01566264236, -74.0078885037, -12.5638793251, 64.5935069551, -0.500332628385};
test_label[2355] = '{64.5935069551};
test_output[2355] = '{20.0588811427};
############ END DEBUG ############*/
test_input[18848:18855] = '{32'h42c44f14, 32'hc212b8f8, 32'hc28e65f0, 32'h4261090c, 32'hc1f9bb6d, 32'hc283b837, 32'h42b0a733, 32'h418ec4a3};
test_label[2356] = '{32'h42b0a733};
test_output[2356] = '{32'h411d3f41};
/*############ DEBUG ############
test_input[18848:18855] = '{98.1544514114, -36.6806322003, -71.1990984288, 56.2588337318, -31.2165173392, -65.8597922365, 88.3265625746, 17.8460142933};
test_label[2356] = '{88.3265625746};
test_output[2356] = '{9.82794276184};
############ END DEBUG ############*/
test_input[18856:18863] = '{32'h4259dd14, 32'h420d0938, 32'h4245a3b1, 32'hc2c3bf9f, 32'hc228c63c, 32'h42a76a4d, 32'hc1d1a839, 32'h41c14182};
test_label[2357] = '{32'hc1d1a839};
test_output[2357] = '{32'h42dbd45b};
/*############ DEBUG ############
test_input[18856:18863] = '{54.4658959288, 35.2590017925, 49.4098561719, -97.8742568151, -42.1935873964, 83.7076189854, -26.2071393517, 24.1569862426};
test_label[2357] = '{-26.2071393517};
test_output[2357] = '{109.914758337};
############ END DEBUG ############*/
test_input[18864:18871] = '{32'h421a6747, 32'h417b184a, 32'hc27e94dc, 32'hc2c723c4, 32'h42afb43f, 32'hc21f74e3, 32'h42853202, 32'h42b450e9};
test_label[2358] = '{32'h421a6747};
test_output[2358] = '{32'h424e9bd3};
/*############ DEBUG ############
test_input[18864:18871] = '{38.6008566565, 15.6934301375, -63.6453701611, -99.5698569337, 87.8520458453, -39.8641471155, 66.5976727977, 90.1580278063};
test_label[2358] = '{38.6008566565};
test_output[2358] = '{51.6521729998};
############ END DEBUG ############*/
test_input[18872:18879] = '{32'h425c1be3, 32'hc1110052, 32'hc243daf1, 32'hc1808d38, 32'h42b6ec81, 32'hc29791b5, 32'hc259e470, 32'hc104b4dd};
test_label[2359] = '{32'hc104b4dd};
test_output[2359] = '{32'h42c7831c};
/*############ DEBUG ############
test_input[18872:18879] = '{55.0272337122, -9.0625783799, -48.9638102527, -16.0689536461, 91.4619179104, -75.7845851502, -54.4730844933, -8.29415583795};
test_label[2359] = '{-8.29415583795};
test_output[2359] = '{99.7560737484};
############ END DEBUG ############*/
test_input[18880:18887] = '{32'hc2ab6704, 32'hc246ea4c, 32'h42995e8e, 32'h41f94780, 32'hc282d748, 32'h42b45281, 32'hc1b3e621, 32'h422d48e7};
test_label[2360] = '{32'hc2ab6704};
test_output[2360] = '{32'h432fdcc3};
/*############ DEBUG ############
test_input[18880:18887] = '{-85.701204393, -49.7288072441, 76.6846755947, 31.1599118766, -65.4204735479, 90.1611426738, -22.4873670716, 43.3211954538};
test_label[2360] = '{-85.701204393};
test_output[2360] = '{175.86234847};
############ END DEBUG ############*/
test_input[18888:18895] = '{32'hc28690ce, 32'h4236ff41, 32'hc21026c8, 32'hc28f3398, 32'hc21057f5, 32'h42319eb1, 32'h41e2809e, 32'h41bfb509};
test_label[2361] = '{32'hc28690ce};
test_output[2361] = '{32'h42e2870e};
/*############ DEBUG ############
test_input[18888:18895] = '{-67.2828250541, 45.7492706007, -36.0378724293, -71.6007710913, -36.0858953318, 44.4049714596, 28.312801636, 23.9633964718};
test_label[2361] = '{-67.2828250541};
test_output[2361] = '{113.263780545};
############ END DEBUG ############*/
test_input[18896:18903] = '{32'h416f6a0d, 32'h42868424, 32'h41130ba7, 32'h421c1242, 32'h4183d821, 32'h42b874a4, 32'h42ad2620, 32'hc2478a62};
test_label[2362] = '{32'h421c1242};
test_output[2362] = '{32'h4254da9b};
/*############ DEBUG ############
test_input[18896:18903] = '{14.9633913225, 67.2580854317, 9.19034459925, 39.0178315511, 16.4805316251, 92.227812604, 86.57446247, -49.8851411892};
test_label[2362] = '{39.0178315511};
test_output[2362] = '{53.2134806744};
############ END DEBUG ############*/
test_input[18904:18911] = '{32'h4194903c, 32'hc2226880, 32'hc1f9289e, 32'h425365c5, 32'hc22c4851, 32'hc2bea697, 32'hc25c37d9, 32'h42089671};
test_label[2363] = '{32'hc2226880};
test_output[2363] = '{32'h42bae722};
/*############ DEBUG ############
test_input[18904:18911] = '{18.5704263175, -40.6020492927, -31.1448331898, 52.849383397, -43.0706230002, -95.3253700648, -55.0545374089, 34.146916767};
test_label[2363] = '{-40.6020492927};
test_output[2363] = '{93.4514326972};
############ END DEBUG ############*/
test_input[18912:18919] = '{32'hc212282a, 32'hc15d0120, 32'hc13010b2, 32'hc094b467, 32'h417b3084, 32'hc25ec5c7, 32'hc2b032fd, 32'hc0c829e4};
test_label[2364] = '{32'hc25ec5c7};
test_output[2364] = '{32'h428ec8f4};
/*############ DEBUG ############
test_input[18912:18919] = '{-36.5392234346, -13.8127742994, -11.0040758065, -4.64702186417, 15.6993450591, -55.6931418611, -88.0995873802, -6.25511364988};
test_label[2364] = '{-55.6931418611};
test_output[2364] = '{71.3924869219};
############ END DEBUG ############*/
test_input[18920:18927] = '{32'hc2a53943, 32'h412a42b9, 32'h426090ff, 32'hc26cb5a8, 32'h41e96a94, 32'h4164d2b3, 32'hc1e6e9da, 32'hc2b7434b};
test_label[2365] = '{32'h412a42b9};
test_output[2365] = '{32'h42360050};
/*############ DEBUG ############
test_input[18920:18927] = '{-82.6118365602, 10.6412897353, 56.1415962512, -59.1773999806, 29.1770398866, 14.3014406186, -28.8641853236, -91.6314286887};
test_label[2365] = '{10.6412897353};
test_output[2365] = '{45.5003065159};
############ END DEBUG ############*/
test_input[18928:18935] = '{32'hc2ac03a1, 32'h423c8c67, 32'h42c17941, 32'h40a53097, 32'h41b60609, 32'hc1cc4623, 32'hc249f355, 32'h42aaaa26};
test_label[2366] = '{32'h42aaaa26};
test_output[2366] = '{32'h413678e6};
/*############ DEBUG ############
test_input[18928:18935] = '{-86.0070868955, 47.1371113752, 96.7368241209, 5.16218150284, 22.7529470171, -25.5342463094, -50.4876290548, 85.3323186976};
test_label[2366] = '{85.3323186976};
test_output[2366] = '{11.4045165684};
############ END DEBUG ############*/
test_input[18936:18943] = '{32'h4263c012, 32'h42576c23, 32'h40ff0410, 32'hc1cd53eb, 32'h42bb33cb, 32'h41997da6, 32'hc2a114a8, 32'h42b9c1a6};
test_label[2367] = '{32'h41997da6};
test_output[2367] = '{32'h42959ef2};
/*############ DEBUG ############
test_input[18936:18943] = '{56.9375678597, 53.8556018861, 7.96924585037, -25.6659761231, 93.6011591364, 19.1863518966, -80.5403467737, 92.8782197582};
test_label[2367] = '{19.1863518966};
test_output[2367] = '{74.810439906};
############ END DEBUG ############*/
test_input[18944:18951] = '{32'hc2bbac44, 32'h4219aec1, 32'hc27101a7, 32'hc29d44bc, 32'h427fcb5d, 32'hc1b2e691, 32'hc25423f4, 32'hc2bd1448};
test_label[2368] = '{32'hc29d44bc};
test_output[2368] = '{32'h430e9535};
/*############ DEBUG ############
test_input[18944:18951] = '{-93.8364573436, 38.4206585926, -60.2516145205, -78.6342460199, 63.9485950673, -22.36258197, -53.0351099411, -94.5396117592};
test_label[2368] = '{-78.6342460199};
test_output[2368] = '{142.582841087};
############ END DEBUG ############*/
test_input[18952:18959] = '{32'h404dfd78, 32'hc2749d42, 32'h42bdc4e8, 32'h419aa2b7, 32'h429c247f, 32'h42c7c513, 32'hc2b356ae, 32'hc213ebdc};
test_label[2369] = '{32'hc2749d42};
test_output[2369] = '{32'h43210b92};
/*############ DEBUG ############
test_input[18952:18959] = '{3.21859550345, -61.1535723185, 94.8845839022, 19.3294513805, 78.0712812982, 99.8849118489, -89.6692987719, -36.9803295265};
test_label[2369] = '{-61.1535723185};
test_output[2369] = '{161.045197322};
############ END DEBUG ############*/
test_input[18960:18967] = '{32'hc2a2fd5d, 32'hc1d0dc65, 32'hc17679be, 32'h41b8a551, 32'h420113ed, 32'h41b92b51, 32'h4195b8bd, 32'hc2158ba1};
test_label[2370] = '{32'hc2a2fd5d};
test_output[2370] = '{32'h42e3876f};
/*############ DEBUG ############
test_input[18960:18967] = '{-81.4948515417, -26.1076141243, -15.4047218937, 23.0807214106, 32.2694570179, 23.1461499855, 18.7152046678, -37.38635647};
test_label[2370] = '{-81.4948515417};
test_output[2370] = '{113.764521113};
############ END DEBUG ############*/
test_input[18968:18975] = '{32'h42a9bbae, 32'hc2bd56b3, 32'hbf398f2c, 32'hc0921d7d, 32'h4290d351, 32'h42a5b024, 32'hc2a8841a, 32'hc2b4032c};
test_label[2371] = '{32'hbf398f2c};
test_output[2371] = '{32'h42ab6e6d};
/*############ DEBUG ############
test_input[18968:18975] = '{84.8665644133, -94.6693373954, -0.724840872605, -4.56609981676, 72.4127305318, 82.8440215147, -84.2580108537, -90.0061957411};
test_label[2371] = '{-0.724840872605};
test_output[2371] = '{85.7156760899};
############ END DEBUG ############*/
test_input[18976:18983] = '{32'hc27033a1, 32'hc28054c4, 32'h411c2a08, 32'h3ff66fca, 32'hc2b0dd27, 32'hc1cbb705, 32'hc23e6378, 32'h419718c0};
test_label[2372] = '{32'hc1cbb705};
test_output[2372] = '{32'h423167ff};
/*############ DEBUG ############
test_input[18976:18983] = '{-60.0504182186, -64.1655571917, 9.76026191106, 1.92528656227, -88.4319383111, -25.4643642238, -47.5971356479, 18.8870848926};
test_label[2372] = '{-25.4643642238};
test_output[2372] = '{44.3515578639};
############ END DEBUG ############*/
test_input[18984:18991] = '{32'h4268ad63, 32'h42473e52, 32'hc294fc64, 32'hc2b495a4, 32'hc23901b7, 32'hc2665d90, 32'h4267fd10, 32'h42a751d7};
test_label[2373] = '{32'hc2665d90};
test_output[2373] = '{32'h430d404f};
/*############ DEBUG ############
test_input[18984:18991] = '{58.1693230558, 49.8108586521, -74.4929539646, -90.2922691683, -46.2516755799, -57.5913680497, 57.9971329988, 83.6598407053};
test_label[2373] = '{-57.5913680497};
test_output[2373] = '{141.251208755};
############ END DEBUG ############*/
test_input[18992:18999] = '{32'hc2720144, 32'hc2812cd1, 32'hc2c12cac, 32'h425f3b9d, 32'h42b5895c, 32'h42b235ba, 32'hc1c649f2, 32'h41e1cd3a};
test_label[2374] = '{32'h425f3b9d};
test_output[2374] = '{32'h420c88cf};
/*############ DEBUG ############
test_input[18992:18999] = '{-60.5012378034, -64.5875335735, -96.5872526357, 55.8082155145, 90.7682815579, 89.1049344919, -24.786105437, 28.2252085739};
test_label[2374] = '{55.8082155145};
test_output[2374] = '{35.1336021511};
############ END DEBUG ############*/
test_input[19000:19007] = '{32'h424a15e8, 32'hc20e5536, 32'hc21d22e3, 32'h42884ba7, 32'h4236ca82, 32'hc126eea5, 32'h4239e6bc, 32'hc299051f};
test_label[2375] = '{32'hc20e5536};
test_output[2375] = '{32'h42cf7642};
/*############ DEBUG ############
test_input[19000:19007] = '{50.5213937067, -35.5832123198, -39.2840698244, 68.1477561814, 45.6977605396, -10.4332632201, 46.4753273057, -76.5100042326};
test_label[2375] = '{-35.5832123198};
test_output[2375] = '{103.730968524};
############ END DEBUG ############*/
test_input[19008:19015] = '{32'hc22ddb32, 32'h4193b571, 32'h4181e675, 32'h429c804c, 32'h42abebe0, 32'hc2c183fe, 32'hc05acf66, 32'hc2a39883};
test_label[2376] = '{32'hc05acf66};
test_output[2376] = '{32'h42b2c296};
/*############ DEBUG ############
test_input[19008:19015] = '{-43.4640571424, 18.4635934846, 16.2375281336, 78.2505820077, 85.960693278, -96.7577942983, -3.41890857535, -81.7978774331};
test_label[2376] = '{-3.41890857535};
test_output[2376] = '{89.3800500245};
############ END DEBUG ############*/
test_input[19016:19023] = '{32'hc294f4a7, 32'h4208d81c, 32'hc1c2255b, 32'hc2b6dd71, 32'hc0852d98, 32'h415a0192, 32'h3f2b19e2, 32'h41d6f953};
test_label[2377] = '{32'h4208d81c};
test_output[2377] = '{32'h3a2a354a};
/*############ DEBUG ############
test_input[19016:19023] = '{-74.477834933, 34.2110440843, -24.2682399224, -91.4325000945, -4.16181576761, 13.6253838344, 0.668363690034, 26.8717398638};
test_label[2377] = '{34.2110440843};
test_output[2377] = '{0.000649292585583};
############ END DEBUG ############*/
test_input[19024:19031] = '{32'h4217e814, 32'hc0ac66eb, 32'hc2c1997a, 32'hc28a1ea7, 32'h4251b694, 32'hc257b6a5, 32'hc29d8e07, 32'h401226c4};
test_label[2378] = '{32'hc257b6a5};
test_output[2378] = '{32'h42d4b69d};
/*############ DEBUG ############
test_input[19024:19031] = '{37.9766378791, -5.38756321768, -96.7997621581, -69.0598664653, 52.4282998755, -53.9283633685, -78.7773946347, 2.28361612738};
test_label[2378] = '{-53.9283633685};
test_output[2378] = '{106.356663773};
############ END DEBUG ############*/
test_input[19032:19039] = '{32'h427e3c79, 32'hc2bbef77, 32'hc20a16a3, 32'hc270bd0e, 32'hc1b60502, 32'hc1d869e8, 32'hc2a95f69, 32'hc288158b};
test_label[2379] = '{32'hc1b60502};
test_output[2379] = '{32'h42ac9f7d};
/*############ DEBUG ############
test_input[19032:19039] = '{63.5590559049, -93.9677072339, -34.5221053584, -60.1846253863, -22.7524457138, -27.0517117431, -84.6863484301, -68.0420723764};
test_label[2379] = '{-22.7524457138};
test_output[2379] = '{86.3115016187};
############ END DEBUG ############*/
test_input[19040:19047] = '{32'h42bf4090, 32'h42c37ec7, 32'hc281dccc, 32'h41a284f3, 32'h42a0341d, 32'hc2bed9d4, 32'h42a8ba5a, 32'hc29a748f};
test_label[2380] = '{32'h42c37ec7};
test_output[2380] = '{32'h3de7d346};
/*############ DEBUG ############
test_input[19040:19047] = '{95.6260967149, 97.7476129454, -64.9312432751, 20.3149174901, 80.1017805839, -95.425445126, 84.3639678845, -77.2276551129};
test_label[2380] = '{97.7476129454};
test_output[2380] = '{0.113195937766};
############ END DEBUG ############*/
test_input[19048:19055] = '{32'h419524ce, 32'h425ff066, 32'hc266b5ce, 32'hc23fc985, 32'hc1b90482, 32'h42986831, 32'hc2922228, 32'h42b8d5c8};
test_label[2381] = '{32'hc23fc985};
test_output[2381] = '{32'h430c5d45};
/*############ DEBUG ############
test_input[19048:19055] = '{18.642970116, 55.9847652406, -57.6775441023, -47.9467958366, -23.1272006201, 76.2034982996, -73.0667098426, 92.4175397738};
test_label[2381] = '{-47.9467958366};
test_output[2381] = '{140.364335701};
############ END DEBUG ############*/
test_input[19056:19063] = '{32'hc237cd2c, 32'hc1dbe9de, 32'h416ecbe0, 32'h424d725a, 32'h4264ceaa, 32'hbffa707c, 32'hc296d47e, 32'h41d04186};
test_label[2382] = '{32'h41d04186};
test_output[2382] = '{32'h41f961c1};
/*############ DEBUG ############
test_input[19056:19063] = '{-45.9503636655, -27.4891921082, 14.9247740869, 51.3616704597, 57.2018219653, -1.95655772639, -75.4150225345, 26.0319940924};
test_label[2382] = '{26.0319940924};
test_output[2382] = '{31.1727320537};
############ END DEBUG ############*/
test_input[19064:19071] = '{32'h427a14c9, 32'hc26af511, 32'h427da084, 32'h422a1f8c, 32'hc23d1d9c, 32'hc1d412bb, 32'h412abf72, 32'h42144112};
test_label[2383] = '{32'hc1d412bb};
test_output[2383] = '{32'h42b485a0};
/*############ DEBUG ############
test_input[19064:19071] = '{62.5202965353, -58.739322347, 63.4067551245, 42.5308070958, -47.2789142028, -26.5091448397, 10.6717392367, 37.0635451001};
test_label[2383] = '{-26.5091448397};
test_output[2383] = '{90.2609868682};
############ END DEBUG ############*/
test_input[19072:19079] = '{32'h4294aba1, 32'h419ff610, 32'hc213b336, 32'h4201d9a3, 32'hc086b321, 32'h42aa2aea, 32'hc0817912, 32'hc1eef403};
test_label[2384] = '{32'hc086b321};
test_output[2384] = '{32'h42b2961f};
/*############ DEBUG ############
test_input[19072:19079] = '{74.3352140753, 19.9951480106, -36.9250106964, 32.4625359721, -4.20936616364, 85.0838193261, -4.04602887999, -29.8691462976};
test_label[2384] = '{-4.20936616364};
test_output[2384] = '{89.2932069649};
############ END DEBUG ############*/
test_input[19080:19087] = '{32'hc278b2ae, 32'h429d150e, 32'hc2662250, 32'h429ae615, 32'hc2ac4f5a, 32'hc27dae2a, 32'h41f4a73b, 32'hc2a12d02};
test_label[2385] = '{32'h429ae615};
test_output[2385] = '{32'h3fb0c964};
/*############ DEBUG ############
test_input[19080:19087] = '{-62.1744919612, 78.5411246584, -57.5335090127, 77.4493827724, -86.1549864774, -63.4200817286, 30.5816552017, -80.5879060349};
test_label[2385] = '{77.4493827724};
test_output[2385] = '{1.38114598942};
############ END DEBUG ############*/
test_input[19088:19095] = '{32'hc1820f24, 32'hc27dcb76, 32'h41b0718d, 32'hc12d35f1, 32'h42b89876, 32'h428f6786, 32'hc2614294, 32'hc26ebb13};
test_label[2386] = '{32'hc1820f24};
test_output[2386] = '{32'h42d91c3f};
/*############ DEBUG ############
test_input[19088:19095] = '{-16.2573931027, -63.4486937167, 22.0554440278, -10.8256696623, 92.2977742865, 71.7021970186, -56.3150183999, -59.6826901709};
test_label[2386] = '{-16.2573931027};
test_output[2386] = '{108.55516739};
############ END DEBUG ############*/
test_input[19096:19103] = '{32'hc2071128, 32'h402cfff9, 32'hc2b28655, 32'hc299da61, 32'hc2aa44f5, 32'hc22b0398, 32'h42c32cbe, 32'hc24cbcb2};
test_label[2387] = '{32'hc2b28655};
test_output[2387] = '{32'h433ad989};
/*############ DEBUG ############
test_input[19096:19103] = '{-33.7667523899, 2.70312327988, -89.2623642706, -76.9265178084, -85.1346817202, -42.7535090449, 97.5873867856, -51.1842714584};
test_label[2387] = '{-89.2623642706};
test_output[2387] = '{186.849751056};
############ END DEBUG ############*/
test_input[19104:19111] = '{32'hc2bdfa5b, 32'h428660a9, 32'hc184b17c, 32'hc0f3b029, 32'hc2a5d563, 32'h40aa3267, 32'h42642e00, 32'hc1b36ce2};
test_label[2388] = '{32'hc184b17c};
test_output[2388] = '{32'h42a78d0d};
/*############ DEBUG ############
test_input[19104:19111] = '{-94.9889741072, 67.1887910834, -16.5866623551, -7.61525373651, -82.916770835, 5.31865245359, 57.0449228791, -22.4281645737};
test_label[2388] = '{-16.5866623551};
test_output[2388] = '{83.7754927542};
############ END DEBUG ############*/
test_input[19112:19119] = '{32'hc2b5bed6, 32'h42557ec8, 32'h417fdd85, 32'hc2a52bdc, 32'h42afbd8f, 32'hc26d3164, 32'h42bf4062, 32'h42a58d5b};
test_label[2389] = '{32'h42557ec8};
test_output[2389] = '{32'h4229026d};
/*############ DEBUG ############
test_input[19112:19119] = '{-90.8727299485, 53.3738092264, 15.9915817312, -82.5856595398, 87.8702295951, -59.2982319651, 95.6257459696, 82.7760853541};
test_label[2389] = '{53.3738092264};
test_output[2389] = '{42.2523676503};
############ END DEBUG ############*/
test_input[19120:19127] = '{32'h42345872, 32'h4220c7de, 32'h41353584, 32'h40f74b02, 32'h41c04a1f, 32'h4158665f, 32'hc25ceddc, 32'h421b3608};
test_label[2390] = '{32'h421b3608};
test_output[2390] = '{32'h40c95fcc};
/*############ DEBUG ############
test_input[19120:19127] = '{45.0863731221, 40.1951824228, 11.3255648933, 7.72790599933, 24.0361920144, 13.5249926771, -55.2322862927, 38.8027647245};
test_label[2390] = '{38.8027647245};
test_output[2390] = '{6.29294381234};
############ END DEBUG ############*/
test_input[19128:19135] = '{32'h42b18381, 32'h417b1a89, 32'hc1f73f06, 32'hc2b6a009, 32'h41af9d77, 32'h4159eb4a, 32'hc2a9e07c, 32'hc1ff0486};
test_label[2391] = '{32'hc2a9e07c};
test_output[2391] = '{32'h432db1fe};
/*############ DEBUG ############
test_input[19128:19135] = '{88.7568411418, 15.6939786284, -30.9057722779, -91.3125694827, 21.9518864877, 13.6199432286, -84.9384434779, -31.8772088833};
test_label[2391] = '{-84.9384434779};
test_output[2391] = '{173.69528462};
############ END DEBUG ############*/
test_input[19136:19143] = '{32'hc25e858b, 32'h4290ef70, 32'hc29e2c29, 32'hc29a0906, 32'h411e0543, 32'hc2508c91, 32'hc259323a, 32'h423e76ef};
test_label[2392] = '{32'hc29a0906};
test_output[2392] = '{32'h43157c3b};
/*############ DEBUG ############
test_input[19136:19143] = '{-55.6304135932, 72.4676529224, -79.0862506473, -77.0176228351, 9.87628426533, -52.1372734813, -54.2990474898, 47.6161456722};
test_label[2392] = '{-77.0176228351};
test_output[2392] = '{149.485275757};
############ END DEBUG ############*/
test_input[19144:19151] = '{32'h428b5b14, 32'h424f20d6, 32'h429d0ffc, 32'h42165117, 32'h4220bce1, 32'h4215ae84, 32'h423887eb, 32'h42ba9b2e};
test_label[2393] = '{32'h4220bce1};
test_output[2393] = '{32'h4254797c};
/*############ DEBUG ############
test_input[19144:19151] = '{69.6778838044, 51.7820656999, 78.5312167925, 37.5791887072, 40.1844506202, 37.420426751, 46.1327307469, 93.3030880293};
test_label[2393] = '{40.1844506202};
test_output[2393] = '{53.1186377934};
############ END DEBUG ############*/
test_input[19152:19159] = '{32'hc2152745, 32'hc2a9c1dc, 32'hc248b97a, 32'hc2478bda, 32'h4204af5f, 32'hc00a91dd, 32'hc2677522, 32'hc2a5b8fa};
test_label[2394] = '{32'hc2a5b8fa};
test_output[2394] = '{32'h42e810aa};
/*############ DEBUG ############
test_input[19152:19159] = '{-37.2883509825, -84.8786304723, -50.1811277058, -49.8865753887, 33.171259095, -2.16515279439, -57.8643888738, -82.8612843134};
test_label[2394] = '{-82.8612843134};
test_output[2394] = '{116.032543408};
############ END DEBUG ############*/
test_input[19160:19167] = '{32'h422be529, 32'h4274ed02, 32'hc10123bd, 32'hc0ef7f1f, 32'h4113a13a, 32'hc10df8f0, 32'h42113d78, 32'hc2b2f058};
test_label[2395] = '{32'h4113a13a};
test_output[2395] = '{32'h425004b3};
/*############ DEBUG ############
test_input[19160:19167] = '{42.9737879547, 61.2314524752, -8.07122542703, -7.48426761788, 9.22686212836, -8.87327551276, 36.3100289375, -89.4694251319};
test_label[2395] = '{9.22686212836};
test_output[2395] = '{52.0045903586};
############ END DEBUG ############*/
test_input[19168:19175] = '{32'h41ca7ade, 32'hc2c5838d, 32'hc218b4f5, 32'h41fa98d3, 32'h42c36d3a, 32'h42baae21, 32'hc27645b8, 32'h41c4c405};
test_label[2396] = '{32'h41fa98d3};
test_output[2396] = '{32'h4284cd6f};
/*############ DEBUG ############
test_input[19168:19175] = '{25.3099930151, -98.7569341508, -38.1767144103, 31.3246215123, 97.7133293217, 93.3400947267, -61.5680865121, 24.5957127846};
test_label[2396] = '{31.3246215123};
test_output[2396] = '{66.4012393457};
############ END DEBUG ############*/
test_input[19176:19183] = '{32'h42c5b751, 32'h42c5ab65, 32'h4274d6a1, 32'h42bf5faa, 32'h428280c4, 32'h42253fe2, 32'h429e8f1c, 32'h422b68e4};
test_label[2397] = '{32'h42c5ab65};
test_output[2397] = '{32'h3f39d1ae};
/*############ DEBUG ############
test_input[19176:19183] = '{98.8580386097, 98.8347548479, 61.2096000552, 95.6868437186, 65.2514978131, 41.3123840498, 79.2795121735, 42.852433177};
test_label[2397] = '{98.8347548479};
test_output[2397] = '{0.725855716629};
############ END DEBUG ############*/
test_input[19184:19191] = '{32'hc2a642b8, 32'hc21035b1, 32'h42954b8b, 32'hc2b09ea9, 32'h41fdf702, 32'h41b4e8ba, 32'hc2550356, 32'hc2347106};
test_label[2398] = '{32'h41b4e8ba};
test_output[2398] = '{32'h425022b8};
/*############ DEBUG ############
test_input[19184:19191] = '{-83.1303068502, -36.0524324655, 74.6475420413, -88.309883581, 31.7456084149, 22.613636006, -53.2532575731, -45.1103744168};
test_label[2398] = '{22.613636006};
test_output[2398] = '{52.0339060353};
############ END DEBUG ############*/
test_input[19192:19199] = '{32'h41f1e2c0, 32'hc2c05a99, 32'hc2bfbb1d, 32'h42725c30, 32'hc1eaa2c3, 32'h4225bea2, 32'hc28bc999, 32'hc26fe862};
test_label[2399] = '{32'hc1eaa2c3};
test_output[2399] = '{32'h42b3d6c9};
/*############ DEBUG ############
test_input[19192:19199] = '{30.2357175763, -96.176945474, -95.8654554483, 60.5900269364, -29.32947301, 41.4361636832, -69.8937486298, -59.9769377911};
test_label[2399] = '{-29.32947301};
test_output[2399] = '{89.9194999512};
############ END DEBUG ############*/
test_input[19200:19207] = '{32'hc2a7a952, 32'hc1ea6c67, 32'h424d3fa0, 32'hc1f51ad2, 32'hc2b24fbf, 32'h42b3e927, 32'hc24f11f9, 32'hc2a5e35d};
test_label[2400] = '{32'hc2a7a952};
test_output[2400] = '{32'h432dc93c};
/*############ DEBUG ############
test_input[19200:19207] = '{-83.8307024956, -29.3029298851, 51.3121352281, -30.6380965667, -89.1557573314, 89.955375824, -51.7675502596, -82.9440656144};
test_label[2400] = '{-83.8307024956};
test_output[2400] = '{173.78607832};
############ END DEBUG ############*/
test_input[19208:19215] = '{32'hc0f90335, 32'h4276dc5b, 32'hc12b93a4, 32'hc29b4b7a, 32'h410361af, 32'h42975c2b, 32'h42b52cd9, 32'hc291b953};
test_label[2401] = '{32'hc29b4b7a};
test_output[2401] = '{32'h43283c2a};
/*############ DEBUG ############
test_input[19208:19215] = '{-7.78164156381, 61.7151922349, -10.7235451888, -77.6474121654, 8.21134834913, 75.6800164406, 90.5875965964, -72.86196118};
test_label[2401] = '{-77.6474121654};
test_output[2401] = '{168.235009097};
############ END DEBUG ############*/
test_input[19216:19223] = '{32'h42a0416e, 32'h42ad7789, 32'h428f9d6c, 32'h425d4302, 32'hc2b603d0, 32'h422d2130, 32'h41c5d3c9, 32'hc24b49c9};
test_label[2402] = '{32'h428f9d6c};
test_output[2402] = '{32'h416ed672};
/*############ DEBUG ############
test_input[19216:19223] = '{80.1277917566, 86.7334697283, 71.8074666447, 55.3154381344, -91.0074428745, 43.2824087801, 24.7284112327, -50.822055801};
test_label[2402] = '{71.8074666447};
test_output[2402] = '{14.9273551644};
############ END DEBUG ############*/
test_input[19224:19231] = '{32'h42bd483d, 32'h429f8198, 32'hc288f750, 32'h42885e82, 32'hc1c51e16, 32'h4262d8cb, 32'hc298adcf, 32'hc22ca15e};
test_label[2403] = '{32'h42885e82};
test_output[2403] = '{32'h41d3a6ed};
/*############ DEBUG ############
test_input[19224:19231] = '{94.6410921503, 79.7531122896, -68.4830347476, 68.184584914, -24.6396901828, 56.7117120324, -76.3394724465, -43.1575853028};
test_label[2403] = '{68.184584914};
test_output[2403] = '{26.4565075784};
############ END DEBUG ############*/
test_input[19232:19239] = '{32'hc11cae06, 32'hc2c6c376, 32'hc2c290d5, 32'h41839a48, 32'h42ab6bd7, 32'hc252d863, 32'h42b831f2, 32'hc161764d};
test_label[2404] = '{32'h42ab6bd7};
test_output[2404] = '{32'h40cc6f6d};
/*############ DEBUG ############
test_input[19232:19239] = '{-9.79248618069, -99.3817560582, -97.2828747749, 16.4503317931, 85.7106272486, -52.7113152209, 92.0975472073, -14.0913820614};
test_label[2404] = '{85.7106272486};
test_output[2404] = '{6.38860197659};
############ END DEBUG ############*/
test_input[19240:19247] = '{32'hc2b9da84, 32'h415dd5dc, 32'h419bdfb7, 32'h42174526, 32'h42bfc8ca, 32'hc0b3e6e8, 32'hc1f3bca4, 32'h413b6ce1};
test_label[2405] = '{32'h413b6ce1};
test_output[2405] = '{32'h42a85b2e};
/*############ DEBUG ############
test_input[19240:19247] = '{-92.9267919232, 13.8647116411, 19.4842365538, 37.8175295924, 95.8921674204, -5.6219368027, -30.467110199, 11.7140821133};
test_label[2405] = '{11.7140821133};
test_output[2405] = '{84.178085307};
############ END DEBUG ############*/
test_input[19248:19255] = '{32'h42987bcf, 32'h421b5f17, 32'h4114543f, 32'hc2bcb6ad, 32'hc28a7ad4, 32'h421b159f, 32'hc21abfcf, 32'h4283bd9d};
test_label[2406] = '{32'hc2bcb6ad};
test_output[2406] = '{32'h432a9940};
/*############ DEBUG ############
test_input[19248:19255] = '{76.2418117163, 38.8428607996, 9.27056802739, -94.3567874327, -69.2398958147, 38.771115133, -38.6873139967, 65.8703378353};
test_label[2406] = '{-94.3567874327};
test_output[2406] = '{170.598630462};
############ END DEBUG ############*/
test_input[19256:19263] = '{32'hc2334911, 32'h3df92639, 32'hc1a50e8b, 32'hc2908e46, 32'hc2a9cfcc, 32'h4135940e, 32'hc1f8b3ff, 32'h42bb8106};
test_label[2407] = '{32'h42bb8106};
test_output[2407] = '{32'h80000000};
/*############ DEBUG ############
test_input[19256:19263] = '{-44.8213538853, 0.121654933964, -20.632101771, -72.2778785051, -84.9058544223, 11.3486457099, -31.0878896041, 93.7519986163};
test_label[2407] = '{93.7519986163};
test_output[2407] = '{-0.0};
############ END DEBUG ############*/
test_input[19264:19271] = '{32'h42673233, 32'h424fd028, 32'hc28b9fe2, 32'hc2b36ad5, 32'hc0dcd301, 32'h41161b13, 32'h42bd9101, 32'h41f1e94f};
test_label[2408] = '{32'hc0dcd301};
test_output[2408] = '{32'h42cb5e32};
/*############ DEBUG ############
test_input[19264:19271] = '{57.7990225534, 51.9532780117, -69.8122706409, -89.7086594372, -6.90075738725, 9.38160982851, 94.7832141043, 30.2389198059};
test_label[2408] = '{-6.90075738725};
test_output[2408] = '{101.683971492};
############ END DEBUG ############*/
test_input[19272:19279] = '{32'h41d99351, 32'hbf917c79, 32'hc26bb0e7, 32'h42888ac2, 32'h420813ef, 32'h42b3aaed, 32'hc1efae40, 32'h42201b0a};
test_label[2409] = '{32'hbf917c79};
test_output[2409] = '{32'h42b5f0df};
/*############ DEBUG ############
test_input[19272:19279] = '{27.1969311217, -1.13661105971, -58.9227556445, 68.2710123686, 34.0194669234, 89.833837177, -29.9600830849, 40.0264066822};
test_label[2409] = '{-1.13661105971};
test_output[2409] = '{90.9704482371};
############ END DEBUG ############*/
test_input[19280:19287] = '{32'hc1b2b75c, 32'hc2b9d7e5, 32'hc1fa4d33, 32'h42c3d3eb, 32'hc2097d45, 32'hc2a803b9, 32'hc2b0e1d3, 32'h42c52630};
test_label[2410] = '{32'hc1b2b75c};
test_output[2410] = '{32'h42f2a93a};
/*############ DEBUG ############
test_input[19280:19287] = '{-22.3395314103, -92.9216720542, -31.287694732, 97.9138991164, -34.3723335033, -84.0072686126, -88.4410664478, 98.5745876183};
test_label[2410] = '{-22.3395314103};
test_output[2410] = '{121.330521178};
############ END DEBUG ############*/
test_input[19288:19295] = '{32'hc1a348c5, 32'h4289b222, 32'h41faa66f, 32'h4282f6a8, 32'h4244a2f3, 32'hc2525e3c, 32'hc2b5d37b, 32'hc2b64e72};
test_label[2411] = '{32'hc1a348c5};
test_output[2411] = '{32'h42b295b4};
/*############ DEBUG ############
test_input[19288:19295] = '{-20.4105315336, 68.8479190026, 31.3312666399, 65.4817502018, 49.1591312052, -52.5920242225, -90.9130476731, -91.1532102847};
test_label[2411] = '{-20.4105315336};
test_output[2411] = '{89.2923896787};
############ END DEBUG ############*/
test_input[19296:19303] = '{32'hc18c10b7, 32'hc20acff6, 32'hc2393b58, 32'h41b6bf2d, 32'h42bbb817, 32'hc286aa2d, 32'hc187c81d, 32'h42a3f104};
test_label[2412] = '{32'hc2393b58};
test_output[2412] = '{32'h430c2ae2};
/*############ DEBUG ############
test_input[19296:19303] = '{-17.5081618354, -34.7030860337, -46.3079546453, 22.8433474397, 93.8595498495, -67.3323765927, -16.9727116601, 81.97073295};
test_label[2412] = '{-46.3079546453};
test_output[2412] = '{140.167511362};
############ END DEBUG ############*/
test_input[19304:19311] = '{32'h40188f48, 32'hc26cd921, 32'h41e76386, 32'h41d0d124, 32'hc11bbde9, 32'hc24128aa, 32'hc2af3c5a, 32'hc27e526c};
test_label[2413] = '{32'h40188f48};
test_output[2413] = '{32'h41d4c804};
/*############ DEBUG ############
test_input[19304:19311] = '{2.38374528304, -59.212041535, 28.9235946367, 26.1021191124, -9.73386447443, -48.2897107555, -87.6178767372, -63.5804901747};
test_label[2413] = '{2.38374528304};
test_output[2413] = '{26.5976634957};
############ END DEBUG ############*/
test_input[19312:19319] = '{32'hc2b106e0, 32'h420d3ca1, 32'h425ea93e, 32'h429bc8a4, 32'hc19bb8a4, 32'hc1b6882e, 32'h3fe45f6a, 32'hc2517c45};
test_label[2414] = '{32'h429bc8a4};
test_output[2414] = '{32'h2f748480};
/*############ DEBUG ############
test_input[19312:19319] = '{-88.5134253867, 35.3092060853, 55.6652743454, 77.8918746688, -19.4651567399, -22.816494594, 1.78416180493, -52.3713582925};
test_label[2414] = '{77.8918746688};
test_output[2414] = '{2.2238744182e-10};
############ END DEBUG ############*/
test_input[19320:19327] = '{32'hc2acd63c, 32'h420a8408, 32'h42bfb16a, 32'hc29797a6, 32'h4246f74a, 32'hc1fb9c7c, 32'hc0f85d14, 32'hc26936c3};
test_label[2415] = '{32'h4246f74a};
test_output[2415] = '{32'h42386b89};
/*############ DEBUG ############
test_input[19320:19327] = '{-86.4184289981, 34.6289363023, 95.8465085811, -75.7961852315, 49.7414934244, -31.4514076089, -7.76136221361, -58.3034781439};
test_label[2415] = '{49.7414934244};
test_output[2415] = '{46.1050151566};
############ END DEBUG ############*/
test_input[19328:19335] = '{32'hc2376cef, 32'h41f0897c, 32'h42813681, 32'h422df098, 32'hc18163e5, 32'h42a7b922, 32'hc19b9c5a, 32'h42c65f49};
test_label[2416] = '{32'h422df098};
test_output[2416] = '{32'h425ecdfa};
/*############ DEBUG ############
test_input[19328:19335] = '{-45.8563802115, 30.0671315292, 64.6064533441, 43.4849549382, -16.1737762079, 83.8615857589, -19.4513430932, 99.1861031216};
test_label[2416] = '{43.4849549382};
test_output[2416] = '{55.7011484046};
############ END DEBUG ############*/
test_input[19336:19343] = '{32'hc2a91e4a, 32'hc202c370, 32'h4223c03b, 32'hc216831a, 32'h40cb25cc, 32'h4268133a, 32'hc246f216, 32'h42a1a091};
test_label[2417] = '{32'hc2a91e4a};
test_output[2417] = '{32'h43255f6e};
/*############ DEBUG ############
test_input[19336:19343] = '{-84.5591563653, -32.6908577073, 40.9377242509, -37.6280282694, 6.34836392386, 58.0187776877, -49.7364113814, 80.8136090682};
test_label[2417] = '{-84.5591563653};
test_output[2417] = '{165.372765434};
############ END DEBUG ############*/
test_input[19344:19351] = '{32'h428ee560, 32'h426174e5, 32'h427b15ac, 32'hc1b5872c, 32'h42512c54, 32'hc1a350fa, 32'hc1a62476, 32'h4274241d};
test_label[2418] = '{32'hc1b5872c};
test_output[2418] = '{32'h42bc4745};
/*############ DEBUG ############
test_input[19344:19351] = '{71.4479977824, 56.3641558325, 62.7711626523, -22.6910016528, 52.293288877, -20.4145388791, -20.7678028865, 61.0352654328};
test_label[2418] = '{-22.6910016528};
test_output[2418] = '{94.1392002385};
############ END DEBUG ############*/
test_input[19352:19359] = '{32'h42a1942f, 32'hc1ceda85, 32'hc2733168, 32'hc1693535, 32'h40a5a9b2, 32'h424de06f, 32'h427fd533, 32'hc2b60885};
test_label[2419] = '{32'hc1ceda85};
test_output[2419] = '{32'h42d54ad1};
/*############ DEBUG ############
test_input[19352:19359] = '{80.7894230887, -25.8566997805, -60.7982472641, -14.5754898647, 5.17696492853, 51.4691719739, 63.9582034847, -91.0166384698};
test_label[2419] = '{-25.8566997805};
test_output[2419] = '{106.646122918};
############ END DEBUG ############*/
test_input[19360:19367] = '{32'hc170d815, 32'h41fccaaa, 32'hc2119556, 32'h4225ea3e, 32'h41a244b1, 32'h42c1433b, 32'h41eb1bab, 32'hbf9f04f7};
test_label[2420] = '{32'hc170d815};
test_output[2420] = '{32'h42df5e3e};
/*############ DEBUG ############
test_input[19360:19367] = '{-15.0527540615, 31.598957111, -36.3958353264, 41.4787521474, 20.2835399288, 96.6313105359, 29.3885106787, -1.24233906204};
test_label[2420] = '{-15.0527540615};
test_output[2420] = '{111.684064597};
############ END DEBUG ############*/
test_input[19368:19375] = '{32'hc20be6cd, 32'h427671e3, 32'h4292f4f0, 32'hc1294cf5, 32'h429d03a5, 32'hc283e10b, 32'h4203718e, 32'hc1c1d652};
test_label[2421] = '{32'h4292f4f0};
test_output[2421] = '{32'h40a120c9};
/*############ DEBUG ############
test_input[19368:19375] = '{-34.9753916999, 61.6112163715, 73.4783917491, -10.5812885166, 78.5071180382, -65.9395351358, 32.8608913951, -24.2296484567};
test_label[2421] = '{73.4783917491};
test_output[2421] = '{5.03525213973};
############ END DEBUG ############*/
test_input[19376:19383] = '{32'h4256bfb4, 32'hc262650c, 32'hc1c1ad81, 32'h40a2d5ac, 32'h40fa652a, 32'hc29225d9, 32'hc2a5cc2e, 32'hc2804e52};
test_label[2422] = '{32'h4256bfb4};
test_output[2422] = '{32'h80000000};
/*############ DEBUG ############
test_input[19376:19383] = '{53.6872110889, -56.5986797424, -24.2097194147, 5.08858319448, 7.82484913839, -73.0739244451, -82.8987856445, -64.1529697416};
test_label[2422] = '{53.6872110889};
test_output[2422] = '{-0.0};
############ END DEBUG ############*/
test_input[19384:19391] = '{32'h41a27177, 32'hc2a291b5, 32'hc1ad19f9, 32'hc1b8b9db, 32'hc1c596d1, 32'hc2a5ec09, 32'h426bece6, 32'hc26eda1a};
test_label[2423] = '{32'h426bece6};
test_output[2423] = '{32'h80000000};
/*############ DEBUG ############
test_input[19384:19391] = '{20.3054028862, -81.2845849841, -21.6376817851, -23.0907491363, -24.6986405918, -82.9610094382, 58.9813455814, -59.7129887052};
test_label[2423] = '{58.9813455814};
test_output[2423] = '{-0.0};
############ END DEBUG ############*/
test_input[19392:19399] = '{32'hc276da45, 32'hc0842f25, 32'h423f6a9c, 32'h4178be90, 32'hc2bfbd4a, 32'hc2ae5039, 32'hc22fca30, 32'h413acc17};
test_label[2424] = '{32'h423f6a9c};
test_output[2424] = '{32'h282c0000};
/*############ DEBUG ############
test_input[19392:19399] = '{-61.7131530476, -4.13075476291, 47.8541125636, 15.546523843, -95.8697047126, -87.1566833453, -43.9474485076, 11.6748270773};
test_label[2424] = '{47.8541125636};
test_output[2424] = '{9.54791801178e-15};
############ END DEBUG ############*/
test_input[19400:19407] = '{32'h41fb4db5, 32'hc2bf391f, 32'hc21f2294, 32'hc2242c69, 32'hc2453675, 32'hc291139a, 32'h41799688, 32'hc0c4200e};
test_label[2425] = '{32'hc2bf391f};
test_output[2425] = '{32'h42fe0c8c};
/*############ DEBUG ############
test_input[19400:19407] = '{31.4129422159, -95.6115610578, -39.7837682632, -41.0433696098, -49.3031797302, -72.5382877438, 15.5992506019, -6.12891316163};
test_label[2425] = '{-95.6115610578};
test_output[2425] = '{127.024503409};
############ END DEBUG ############*/
test_input[19408:19415] = '{32'hc18645af, 32'hc1faabf0, 32'h42bcc4d0, 32'hc2951054, 32'hc2c149a3, 32'hc2188fe7, 32'h428507f4, 32'hc1d91b25};
test_label[2426] = '{32'hc2951054};
test_output[2426] = '{32'h4328ea92};
/*############ DEBUG ############
test_input[19408:19415] = '{-16.78402484, -31.3339537085, 94.3844024993, -74.5318907502, -96.6438234609, -38.1405302421, 66.5155355342, -27.138254258};
test_label[2426] = '{-74.5318907502};
test_output[2426] = '{168.91629325};
############ END DEBUG ############*/
test_input[19416:19423] = '{32'hc1bbc0c7, 32'h42843c7b, 32'h42684cc0, 32'hc18a95bf, 32'h42889422, 32'h415fa07e, 32'hc2b679d0, 32'hc1c6355b};
test_label[2427] = '{32'hc18a95bf};
test_output[2427] = '{32'h42ab70e1};
/*############ DEBUG ############
test_input[19416:19423] = '{-23.4691302442, 66.118129721, 58.0749517313, -17.3231174083, 68.2893234061, 13.976682307, -91.2379116916, -24.7760534217};
test_label[2427] = '{-17.3231174083};
test_output[2427] = '{85.7204680126};
############ END DEBUG ############*/
test_input[19424:19431] = '{32'hc2b0ac41, 32'h429971e8, 32'hc17ef137, 32'h41de5d83, 32'h428981e7, 32'hbe991d6c, 32'h4115f658, 32'h42a770fb};
test_label[2428] = '{32'hbe991d6c};
test_output[2428] = '{32'h42a80a90};
/*############ DEBUG ############
test_input[19424:19431] = '{-88.3364314587, 76.7224737724, -15.9338901395, 27.7956601299, 68.7537123934, -0.299052581695, 9.37264214728, 83.72066158};
test_label[2428] = '{-0.299052581695};
test_output[2428] = '{84.0206275965};
############ END DEBUG ############*/
test_input[19432:19439] = '{32'hc266b11e, 32'hc29c639a, 32'hc1e67e71, 32'hc2b487a5, 32'hc2a8b519, 32'h4286ca40, 32'h4128487e, 32'h41d8fefe};
test_label[2429] = '{32'hc266b11e};
test_output[2429] = '{32'h42fa22cf};
/*############ DEBUG ############
test_input[19432:19439] = '{-57.6729676507, -78.194533164, -28.8117387518, -90.2649327646, -84.35370744, 67.3950181422, 10.5176979781, 27.1245083265};
test_label[2429] = '{-57.6729676507};
test_output[2429] = '{125.067985793};
############ END DEBUG ############*/
test_input[19440:19447] = '{32'h41d18f5b, 32'h42b3ab5f, 32'h40b6d12f, 32'hc0dd3a1e, 32'hc2306946, 32'h42077a04, 32'h418a08fe, 32'hc2afab4c};
test_label[2430] = '{32'h40b6d12f};
test_output[2430] = '{32'h42a83e4d};
/*############ DEBUG ############
test_input[19440:19447] = '{26.1949979897, 89.8347129348, 5.71303503795, -6.91334455369, -44.1028043247, 33.8691542611, 17.2543905484, -87.8345613384};
test_label[2430] = '{5.71303503795};
test_output[2430] = '{84.1216778969};
############ END DEBUG ############*/
test_input[19448:19455] = '{32'h41f24581, 32'h427fc984, 32'h427a0a87, 32'hc2526e0f, 32'hc22381df, 32'hc211f992, 32'h41d7f0c6, 32'hc1959188};
test_label[2431] = '{32'hc22381df};
test_output[2431] = '{32'h42d212e8};
/*############ DEBUG ############
test_input[19448:19455] = '{30.2839376044, 63.9467943144, 62.5102808977, -52.607477815, -40.8768287578, -36.493720635, 26.9925653539, -18.6960604993};
test_label[2431] = '{-40.8768287578};
test_output[2431] = '{105.036922544};
############ END DEBUG ############*/
test_input[19456:19463] = '{32'hc238ab95, 32'hc1519890, 32'hc12ef38c, 32'hc29709d5, 32'h423d4369, 32'h4290b634, 32'hc29c3fe2, 32'h4160c8a1};
test_label[2432] = '{32'h4160c8a1};
test_output[2432] = '{32'h42693a40};
/*############ DEBUG ############
test_input[19456:19463] = '{-46.1675605346, -13.0997466069, -10.9344600621, -75.5192024633, 47.3158292701, 72.3558677086, -78.124768219, 14.0489819767};
test_label[2432] = '{14.0489819767};
test_output[2432] = '{58.3068857318};
############ END DEBUG ############*/
test_input[19464:19471] = '{32'h41fa65b7, 32'hc1e67508, 32'hc29f6400, 32'hc2bbbbab, 32'h422fa158, 32'h422cc966, 32'hc25f076f, 32'h4088a99d};
test_label[2433] = '{32'hc29f6400};
test_output[2433] = '{32'h42f80143};
/*############ DEBUG ############
test_input[19464:19471] = '{31.2996656863, -28.8071437468, -79.695313503, -93.8665377997, 43.9075640535, 43.1966776054, -55.7572583379, 4.27070493262};
test_label[2433] = '{-79.695313503};
test_output[2433] = '{124.002466714};
############ END DEBUG ############*/
test_input[19472:19479] = '{32'h42bf0181, 32'h41ab622e, 32'h426dbf57, 32'hc26c4042, 32'h426809d3, 32'h411bbd48, 32'h429095c3, 32'h4144753c};
test_label[2434] = '{32'h426dbf57};
test_output[2434] = '{32'h421043aa};
/*############ DEBUG ############
test_input[19472:19479] = '{95.5029342557, 21.4229385121, 59.4368542794, -59.0627513655, 58.009592332, 9.73371081274, 72.2925059779, 12.2786220539};
test_label[2434] = '{59.4368542794};
test_output[2434] = '{36.0660799764};
############ END DEBUG ############*/
test_input[19480:19487] = '{32'hc2856bd9, 32'hc0994d04, 32'h421e1596, 32'hc2a9f281, 32'h42742f25, 32'hc245346a, 32'h42960dae, 32'h42afba3c};
test_label[2435] = '{32'h42afba3c};
test_output[2435] = '{32'h36328a01};
/*############ DEBUG ############
test_input[19480:19487] = '{-66.7106390244, -4.79065147478, 39.5210815853, -84.9736380862, 61.0460388902, -49.3011872744, 75.0267184875, 87.8637371753};
test_label[2435] = '{87.8637371753};
test_output[2435] = '{2.66043964094e-06};
############ END DEBUG ############*/
test_input[19488:19495] = '{32'h428d94b8, 32'hc0c292bc, 32'hc13e3358, 32'hc2a01e63, 32'h40252271, 32'hc216e380, 32'h4028e420, 32'h4211b197};
test_label[2436] = '{32'h4211b197};
test_output[2436] = '{32'h420977d9};
/*############ DEBUG ############
test_input[19488:19495] = '{70.7904643688, -6.08041180713, -11.887534945, -80.0593511816, 2.58022714344, -37.7221691078, 2.63892373352, 36.4234270984};
test_label[2436] = '{36.4234270984};
test_output[2436] = '{34.3670372704};
############ END DEBUG ############*/
test_input[19496:19503] = '{32'hc23d87c5, 32'hc0bd4b34, 32'hc2749ef1, 32'h4227c160, 32'hbfb1a5d4, 32'hc28e8938, 32'h4299e835, 32'hc2c3ef7b};
test_label[2437] = '{32'hc23d87c5};
test_output[2437] = '{32'h42f8ac18};
/*############ DEBUG ############
test_input[19496:19503] = '{-47.3825870383, -5.91543021126, -61.1552174229, 41.9388420883, -1.38787317229, -71.2680016552, 76.9535327212, -97.967736771};
test_label[2437] = '{-47.3825870383};
test_output[2437] = '{124.336119759};
############ END DEBUG ############*/
test_input[19504:19511] = '{32'h42c110b1, 32'h41c030ce, 32'h41953aee, 32'hc20f6f8c, 32'hc0e1f489, 32'hc2ae3162, 32'h40b6e915, 32'hc24116d3};
test_label[2438] = '{32'h40b6e915};
test_output[2438] = '{32'h42b5a220};
/*############ DEBUG ############
test_input[19504:19511] = '{96.5326003313, 24.0238306071, 18.6537745503, -35.8589310097, -7.06110033488, -87.0964525571, 5.71595260666, -48.2722888933};
test_label[2438] = '{5.71595260666};
test_output[2438] = '{90.8166477246};
############ END DEBUG ############*/
test_input[19512:19519] = '{32'hc205f1b1, 32'hc2c33780, 32'hc29ebd9a, 32'h42c2eb3e, 32'hc2c041c7, 32'h42afa308, 32'h4299f099, 32'h42369490};
test_label[2439] = '{32'h4299f099};
test_output[2439] = '{32'h41a3eab9};
/*############ DEBUG ############
test_input[19512:19519] = '{-33.4860263828, -97.6083969052, -79.3703183919, 97.4594583675, -96.1284688197, 87.8184209541, 76.9699135333, 45.64508012};
test_label[2439] = '{76.9699135333};
test_output[2439] = '{20.4896098389};
############ END DEBUG ############*/
test_input[19520:19527] = '{32'hc1d2874f, 32'h423011f6, 32'h42c4b28f, 32'h414e51f2, 32'hc21b6bb3, 32'h3feeea76, 32'h427cb20e, 32'hc1091f43};
test_label[2440] = '{32'h423011f6};
test_output[2440] = '{32'h42595329};
/*############ DEBUG ############
test_input[19520:19527] = '{-26.316069072, 44.0175402959, 98.3487502167, 12.8950063274, -38.8551744905, 1.86653020138, 63.1738809851, -8.5701321664};
test_label[2440] = '{44.0175402959};
test_output[2440] = '{54.3312099209};
############ END DEBUG ############*/
test_input[19528:19535] = '{32'hc2b05176, 32'hc19c9bd2, 32'h411a900e, 32'hc06fa3e1, 32'h4274820c, 32'h42abdff8, 32'hc28a0782, 32'hc297544c};
test_label[2441] = '{32'h411a900e};
test_output[2441] = '{32'h42988df6};
/*############ DEBUG ############
test_input[19528:19535] = '{-88.1591023811, -19.5760848394, 9.6601696567, -3.74437737805, 61.1270007614, 85.9374372451, -69.0146620474, -75.6646453503};
test_label[2441] = '{9.6601696567};
test_output[2441] = '{76.2772675884};
############ END DEBUG ############*/
test_input[19536:19543] = '{32'hc25b61aa, 32'h4193da36, 32'h41fa4fea, 32'hc28d12d4, 32'hc2993afb, 32'hc2bcc5fc, 32'hc2c42904, 32'hc269823e};
test_label[2442] = '{32'hc269823e};
test_output[2442] = '{32'h42b3551a};
/*############ DEBUG ############
test_input[19536:19543] = '{-54.8453769035, 18.4815491324, 31.2890214607, -70.5367707031, -76.6151962012, -94.3866865225, -98.0801120107, -58.3771909167};
test_label[2442] = '{-58.3771909167};
test_output[2442] = '{89.6662151176};
############ END DEBUG ############*/
test_input[19544:19551] = '{32'h42bccbd9, 32'hc2a79c86, 32'h428990ab, 32'h41b8df60, 32'hc2b4ac33, 32'hc2886141, 32'hc2a2f58a, 32'h4266c182};
test_label[2443] = '{32'hc2a79c86};
test_output[2443] = '{32'h43323430};
/*############ DEBUG ############
test_input[19544:19551] = '{94.3981392114, -83.8057123022, 68.7825555541, 23.1090702877, -90.3363271055, -68.1899498188, -81.479569566, 57.6889707919};
test_label[2443] = '{-83.8057123022};
test_output[2443] = '{178.203851514};
############ END DEBUG ############*/
test_input[19552:19559] = '{32'h42889fdd, 32'h427afe81, 32'h42b3f08c, 32'hc16b59d0, 32'h4293ae95, 32'hc1f0fe83, 32'h424c10a2, 32'h42bb0f2a};
test_label[2444] = '{32'h4293ae95};
test_output[2444] = '{32'h419dbbc4};
/*############ DEBUG ############
test_input[19552:19559] = '{68.3122356955, 62.7485383304, 89.9698196317, -14.7094268819, 73.8409815273, -30.1242724073, 51.0162422242, 93.5296161454};
test_label[2444] = '{73.8409815273};
test_output[2444] = '{19.7166821965};
############ END DEBUG ############*/
test_input[19560:19567] = '{32'h4296e0df, 32'h42c03711, 32'hc24f271e, 32'h41c29c6a, 32'h4234573e, 32'hc14b8157, 32'hc192b5b2, 32'hc281170a};
test_label[2445] = '{32'h42c03711};
test_output[2445] = '{32'h30913297};
/*############ DEBUG ############
test_input[19560:19567] = '{75.439200647, 96.1075507103, -51.7882001412, 24.3263739523, 45.0851960872, -12.7190767596, -18.3387188747, -64.5449989508};
test_label[2445] = '{96.1075507103};
test_output[2445] = '{1.05645170445e-09};
############ END DEBUG ############*/
test_input[19568:19575] = '{32'hc29e437a, 32'h41e72240, 32'h428cd247, 32'hc2c616e2, 32'h4261691c, 32'hc2c5a317, 32'h41d516df, 32'h41f9ed57};
test_label[2446] = '{32'h428cd247};
test_output[2446] = '{32'h35529f77};
/*############ DEBUG ############
test_input[19568:19575] = '{-79.131791068, 28.8917233913, 70.4106962045, -99.044693859, 56.3526449018, -98.8185359786, 26.6361676329, 31.2408886719};
test_label[2446] = '{70.4106962045};
test_output[2446] = '{7.84631469533e-07};
############ END DEBUG ############*/
test_input[19576:19583] = '{32'hc2ab11a4, 32'h4255fc37, 32'hc249ca88, 32'h42918431, 32'h40db127c, 32'hc298b3a4, 32'hc2aa70de, 32'h42aee2cb};
test_label[2447] = '{32'h42aee2cb};
test_output[2447] = '{32'h34e116f9};
/*############ DEBUG ############
test_input[19576:19583] = '{-85.5344534189, 53.4963039928, -50.4477847058, 72.7581836987, 6.84600641536, -76.350858521, -85.2204432659, 87.4429526097};
test_label[2447] = '{87.4429526097};
test_output[2447] = '{4.19262292511e-07};
############ END DEBUG ############*/
test_input[19584:19591] = '{32'h3f05fa9b, 32'hc0e1d21b, 32'hc16c0ef1, 32'h42a34116, 32'h4254946f, 32'hc2290f0b, 32'h4106fd19, 32'hc29dea2e};
test_label[2448] = '{32'h4106fd19};
test_output[2448] = '{32'h42926173};
/*############ DEBUG ############
test_input[19584:19591] = '{0.523355168334, -7.05689741944, -14.7536477434, 81.6271199223, 53.144953784, -42.2646911776, 8.43679183767, -78.9573810796};
test_label[2448] = '{8.43679183767};
test_output[2448] = '{73.1903280846};
############ END DEBUG ############*/
test_input[19592:19599] = '{32'hc214a5e0, 32'h429db652, 32'hc2b0e699, 32'h42b31ec5, 32'h42164da8, 32'h41833435, 32'hc23b2298, 32'h4237d351};
test_label[2449] = '{32'h42b31ec5};
test_output[2449] = '{32'h37bc5cea};
/*############ DEBUG ############
test_input[19592:19599] = '{-37.1619886149, 78.8560908708, -88.4503839075, 89.5600941443, 37.5758349687, 16.4004916719, -46.7837840594, 45.9563650244};
test_label[2449] = '{89.5600941443};
test_output[2449] = '{2.24546126668e-05};
############ END DEBUG ############*/
test_input[19600:19607] = '{32'h428557fb, 32'hc21eac09, 32'h4198998c, 32'hc235816f, 32'hc2457a67, 32'hc1ebbb9d, 32'hc222ee31, 32'h41a68959};
test_label[2450] = '{32'h4198998c};
test_output[2450] = '{32'h423e632f};
/*############ DEBUG ############
test_input[19600:19607] = '{66.6718337562, -39.6680034112, 19.0749732266, -45.3763998394, -49.3695331552, -29.4666087767, -40.7326086018, 20.817063421};
test_label[2450] = '{19.0749732266};
test_output[2450] = '{47.5968605296};
############ END DEBUG ############*/
test_input[19608:19615] = '{32'hc27f4e10, 32'h420567f3, 32'h41ef8a54, 32'h42b7e74a, 32'h42aa500d, 32'hc2acf0b2, 32'hc269a5ea, 32'h4215f50a};
test_label[2451] = '{32'h4215f50a};
test_output[2451] = '{32'h4259daaf};
/*############ DEBUG ############
test_input[19608:19615] = '{-63.8262315124, 33.35151347, 29.9425437718, 91.9517343263, 85.1563522784, -86.4701045832, -58.4120242493, 37.4892957589};
test_label[2451] = '{37.4892957589};
test_output[2451] = '{54.4635568722};
############ END DEBUG ############*/
test_input[19616:19623] = '{32'h414c8f25, 32'h42425a3a, 32'h42b5091f, 32'hc2508821, 32'h4298e5e2, 32'h41a6653f, 32'h40aa6d82, 32'hc292189c};
test_label[2452] = '{32'h42b5091f};
test_output[2452] = '{32'h35505dfe};
/*############ DEBUG ############
test_input[19616:19623] = '{12.7849473406, 48.588112379, 90.5178112793, -52.1329369186, 76.4489923313, 20.7994361192, 5.32586756376, -73.0480639549};
test_label[2452] = '{90.5178112793};
test_output[2452] = '{7.76228162586e-07};
############ END DEBUG ############*/
test_input[19624:19631] = '{32'h4235fb7c, 32'hc2c72c7e, 32'h427b2ae9, 32'hc242a680, 32'hc166793a, 32'h413ef432, 32'h42526399, 32'h41f1f812};
test_label[2453] = '{32'h427b2ae9};
test_output[2453] = '{32'h381cde12};
/*############ DEBUG ############
test_input[19624:19631] = '{45.4955920259, -99.5868961636, 62.7919053387, -48.6625991009, -14.4045959412, 11.9346181923, 52.5972639012, 30.2461276671};
test_label[2453] = '{62.7919053387};
test_output[2453] = '{3.74001160758e-05};
############ END DEBUG ############*/
test_input[19632:19639] = '{32'h3f671802, 32'h41280340, 32'h42c535a5, 32'h424daaed, 32'h416b0694, 32'hc24179c9, 32'h42c04cf2, 32'h42c5106d};
test_label[2454] = '{32'h416b0694};
test_output[2454] = '{32'h42a93bbe};
/*############ DEBUG ############
test_input[19632:19639] = '{0.90271009928, 10.5007932226, 98.6047713423, 51.4169211041, 14.6891055795, -48.3689308327, 96.1502852451, 98.5320852098};
test_label[2454] = '{14.6891055795};
test_output[2454] = '{84.6166818915};
############ END DEBUG ############*/
test_input[19640:19647] = '{32'h422cd4ff, 32'h41a06fdc, 32'h42b02cbd, 32'h4284ecfd, 32'hc18c6171, 32'hc0464a71, 32'hc074cf84, 32'h410c9771};
test_label[2455] = '{32'h42b02cbd};
test_output[2455] = '{32'h2fdf3c68};
/*############ DEBUG ############
test_input[19640:19647] = '{43.2080055434, 20.0546185326, 88.0873757077, 66.4628651345, -17.5475789669, -3.0982934755, -3.82516571466, 8.78697262271};
test_label[2455] = '{88.0873757077};
test_output[2455] = '{4.06063849294e-10};
############ END DEBUG ############*/
test_input[19648:19655] = '{32'hc2884dc6, 32'hc0e29d57, 32'h429dfc53, 32'h42b84f3b, 32'hc229d558, 32'hc25ba102, 32'hc225247c, 32'hc28abb5e};
test_label[2456] = '{32'hc28abb5e};
test_output[2456] = '{32'h4321854c};
/*############ DEBUG ############
test_input[19648:19655] = '{-68.1519003018, -7.08170661813, 78.992819421, 92.1547454279, -42.4583426834, -54.9072349941, -41.2856284858, -69.3659506784};
test_label[2456] = '{-69.3659506784};
test_output[2456] = '{161.520698029};
############ END DEBUG ############*/
test_input[19656:19663] = '{32'hbf53a818, 32'hc26a6877, 32'hc287adcc, 32'h4250ae11, 32'h40df06ae, 32'hc245efc9, 32'h4294d2c4, 32'hc1b2b4e5};
test_label[2457] = '{32'hc245efc9};
test_output[2457] = '{32'h42f7caa9};
/*############ DEBUG ############
test_input[19656:19663] = '{-0.82678365091, -58.6020175003, -67.8394437209, 52.1699856099, 6.96956559402, -49.4841662533, 74.4116537047, -22.3383278986};
test_label[2457] = '{-49.4841662533};
test_output[2457] = '{123.895819958};
############ END DEBUG ############*/
test_input[19664:19671] = '{32'h42a51897, 32'hc1fb7f64, 32'hc27d5f4b, 32'hc2a8a4ab, 32'h4245f274, 32'h414bc580, 32'h414c0624, 32'h425ae7cc};
test_label[2458] = '{32'hc27d5f4b};
test_output[2458] = '{32'h4311e41e};
/*############ DEBUG ############
test_input[19664:19671] = '{82.5480288708, -31.4372025732, -63.3430598086, -84.3216148232, 49.4867724923, 12.7357177564, 12.7514991101, 54.7263637035};
test_label[2458] = '{-63.3430598086};
test_output[2458] = '{145.891088679};
############ END DEBUG ############*/
test_input[19672:19679] = '{32'h41cf17eb, 32'h4120c186, 32'h42809cd7, 32'h41f55cff, 32'h3f34d063, 32'hc1854579, 32'hc2bb9d2a, 32'hc25f44d1};
test_label[2459] = '{32'h41f55cff};
test_output[2459] = '{32'h42068b2e};
/*############ DEBUG ############
test_input[19672:19679] = '{25.8866789966, 10.0472467033, 64.3063263231, 30.6704076851, 0.706304717863, -16.6589225015, -93.8069610681, -55.8172047916};
test_label[2459] = '{30.6704076851};
test_output[2459] = '{33.635918638};
############ END DEBUG ############*/
test_input[19680:19687] = '{32'h4281d389, 32'hc2a51614, 32'h42a00b37, 32'hc27290ac, 32'hc1a35873, 32'h41e85e16, 32'hc2a74c1e, 32'h41a97dfd};
test_label[2460] = '{32'h41e85e16};
test_output[2460] = '{32'h424be764};
/*############ DEBUG ############
test_input[19680:19687] = '{64.9131583745, -82.543120943, 80.0219071463, -60.6412827079, -20.4181879095, 29.04594013, -83.6486650998, 21.1865177582};
test_label[2460] = '{29.04594013};
test_output[2460] = '{50.9759672907};
############ END DEBUG ############*/
test_input[19688:19695] = '{32'h42b23905, 32'hc2b1fbd9, 32'hc275e2bb, 32'h42a2d352, 32'h42179450, 32'hc2af5036, 32'hc248a835, 32'h4273abfd};
test_label[2461] = '{32'h4273abfd};
test_output[2461] = '{32'h41e18d09};
/*############ DEBUG ############
test_input[19688:19695] = '{89.1113661693, -88.9918888737, -61.471416191, 81.4127367881, 37.894835809, -87.65666008, -50.1642639502, 60.9179555554};
test_label[2461] = '{60.9179555554};
test_output[2461] = '{28.1938639594};
############ END DEBUG ############*/
test_input[19696:19703] = '{32'h4235bd98, 32'hc2c0d89e, 32'h42a2c161, 32'hc28f699b, 32'h41c7cd5e, 32'h42af7320, 32'h417d50e3, 32'h42881064};
test_label[2462] = '{32'h41c7cd5e};
test_output[2462] = '{32'h427b015b};
/*############ DEBUG ############
test_input[19696:19703] = '{45.4351514711, -96.4230771834, 81.3776945901, -71.7062598271, 24.9752767268, 87.7248511309, 15.8322476552, 68.0320128017};
test_label[2462] = '{24.9752767268};
test_output[2462] = '{62.7513245954};
############ END DEBUG ############*/
test_input[19704:19711] = '{32'h41811faa, 32'hc2a7f27e, 32'h420a68af, 32'hc2befa88, 32'hc27819ab, 32'hc290d424, 32'hbf53a776, 32'hc2b970e2};
test_label[2463] = '{32'hc2b970e2};
test_output[2463] = '{32'h42fea53a};
/*############ DEBUG ############
test_input[19704:19711] = '{16.1404602856, -83.9736191516, 34.6022318298, -95.4893165483, -62.0250682603, -72.4143406477, -0.826774005272, -92.7204724914};
test_label[2463] = '{-92.7204724914};
test_output[2463] = '{127.322704331};
############ END DEBUG ############*/
test_input[19712:19719] = '{32'h421eb406, 32'h42066b0c, 32'h41d2e210, 32'h41bc848b, 32'hc2adc2c1, 32'hc2a6a246, 32'h427d2070, 32'h429ab45e};
test_label[2464] = '{32'h427d2070};
test_output[2464] = '{32'h41612136};
/*############ DEBUG ############
test_input[19712:19719] = '{39.6758051022, 33.6045365286, 26.3603829886, 23.5647175436, -86.8803783096, -83.3169428312, 63.2816762933, 77.3522832452};
test_label[2464] = '{63.2816762933};
test_output[2464] = '{14.0706077267};
############ END DEBUG ############*/
test_input[19720:19727] = '{32'h42bbe6a5, 32'h418c78fd, 32'h4279dc7c, 32'h41ec3009, 32'hc1994ee1, 32'hc246feae, 32'hc25661da, 32'h42a89e19};
test_label[2465] = '{32'h42bbe6a5};
test_output[2465] = '{32'h38883bd5};
/*############ DEBUG ############
test_input[19720:19727] = '{93.9504740034, 17.5590765529, 62.4653150339, 29.5234544918, -19.1635141778, -49.7487122234, -53.5955569541, 84.3087876129};
test_label[2465] = '{93.9504740034};
test_output[2465] = '{6.49612986403e-05};
############ END DEBUG ############*/
test_input[19728:19735] = '{32'h427049fa, 32'hc0d4acf9, 32'h3fcb5be6, 32'hc1b0356d, 32'hc1957ea7, 32'hc1cfeeb3, 32'h42975229, 32'h41ad575b};
test_label[2466] = '{32'hc0d4acf9};
test_output[2466] = '{32'h42a49cf9};
/*############ DEBUG ############
test_input[19728:19735] = '{60.0722439886, -6.64611499414, 1.5887419921, -22.0260859427, -18.6868423612, -25.9915527231, 75.6604683036, 21.6676535631};
test_label[2466] = '{-6.64611499414};
test_output[2466] = '{82.3065834676};
############ END DEBUG ############*/
test_input[19736:19743] = '{32'h428965ba, 32'h42935356, 32'h41bf17a2, 32'h42181fc0, 32'hc25f7dff, 32'hc221f69c, 32'hc1fd935d, 32'hc18433a6};
test_label[2467] = '{32'hc18433a6};
test_output[2467] = '{32'h42b463d0};
/*############ DEBUG ############
test_input[19736:19743] = '{68.6986827267, 73.6627693104, 23.8865399741, 38.0310056544, -55.873043226, -40.4908305066, -31.6969540944, -16.5252198953};
test_label[2467] = '{-16.5252198953};
test_output[2467] = '{90.1949492557};
############ END DEBUG ############*/
test_input[19744:19751] = '{32'hc2916585, 32'h4171c073, 32'h428711c1, 32'h41822646, 32'h4247bd8d, 32'h40a8ac9a, 32'hc20799d3, 32'hc29e6c8f};
test_label[2468] = '{32'hc20799d3};
test_output[2468] = '{32'h42cadeaa};
/*############ DEBUG ############
test_input[19744:19751] = '{-72.6982768611, 15.109484635, 67.5346739242, 16.2686879542, 49.9351083541, 5.27106955783, -33.900217166, -79.2120266207};
test_label[2468] = '{-33.900217166};
test_output[2468] = '{101.434891113};
############ END DEBUG ############*/
test_input[19752:19759] = '{32'h3e593835, 32'h408dc836, 32'h401448c2, 32'hc2097371, 32'hc2ab4302, 32'hc224e784, 32'hc247adbe, 32'h41bafa6b};
test_label[2469] = '{32'h401448c2};
test_output[2469] = '{32'h41a87153};
/*############ DEBUG ############
test_input[19752:19759] = '{0.212128472895, 4.43069000882, 2.31694090163, -34.3627370142, -85.6308734901, -41.2260912445, -49.919670628, 23.3722747747};
test_label[2469] = '{2.31694090163};
test_output[2469] = '{21.0553338798};
############ END DEBUG ############*/
test_input[19760:19767] = '{32'h418597e7, 32'h4219d07d, 32'hc129dc29, 32'hc234b1fb, 32'hc103b8dd, 32'h413e050a, 32'hc1bba218, 32'h422ae195};
test_label[2470] = '{32'hc234b1fb};
test_output[2470] = '{32'h42afd0ea};
/*############ DEBUG ############
test_input[19760:19767] = '{16.6991705083, 38.4536012263, -10.6162503439, -45.1738098898, -8.23263306543, 11.8762301064, -23.4541481291, 42.7202958399};
test_label[2470] = '{-45.1738098898};
test_output[2470] = '{87.9080363217};
############ END DEBUG ############*/
test_input[19768:19775] = '{32'h42c553b5, 32'hc238b726, 32'hc2baea7e, 32'hc1a33876, 32'hc188a552, 32'h3ed909bb, 32'h41aacdbe, 32'hc0f08ce2};
test_label[2471] = '{32'h42c553b5};
test_output[2471] = '{32'h80000000};
/*############ DEBUG ############
test_input[19768:19775] = '{98.6634884003, -46.1788547054, -93.4579926307, -20.4025693647, -17.0807220296, 0.423902348519, 21.3504592169, -7.51719752558};
test_label[2471] = '{98.6634884003};
test_output[2471] = '{-0.0};
############ END DEBUG ############*/
test_input[19776:19783] = '{32'hc280dfb5, 32'hc2b81626, 32'h40af7419, 32'hc292d0ee, 32'h41fad39d, 32'hc2737802, 32'h4186948f, 32'hc2b3a35d};
test_label[2472] = '{32'hc2b3a35d};
test_output[2472] = '{32'h42f25844};
/*############ DEBUG ############
test_input[19776:19783] = '{-64.4369307277, -92.0432564183, 5.48292212139, -73.4080649652, 31.3533274925, -60.8671951289, 16.8225382678, -89.8190652828};
test_label[2472] = '{-89.8190652828};
test_output[2472] = '{121.172393264};
############ END DEBUG ############*/
test_input[19784:19791] = '{32'h426c6d19, 32'hc2022bd5, 32'h42c500d0, 32'hc06c4d93, 32'hc2a264be, 32'h41590d54, 32'h42a7403d, 32'hc1c79004};
test_label[2473] = '{32'hc06c4d93};
test_output[2473] = '{32'h42cc633d};
/*############ DEBUG ############
test_input[19784:19791] = '{59.1065392651, -32.5428047627, 98.5015886948, -3.69223481532, -81.1967584564, 13.5657542968, 83.6254680878, -24.9453205778};
test_label[2473] = '{-3.69223481532};
test_output[2473] = '{102.193823856};
############ END DEBUG ############*/
test_input[19792:19799] = '{32'h42001bd5, 32'hc2c3d93c, 32'h42b07886, 32'h4283836c, 32'h42840304, 32'hc2215b60, 32'h4190e8ff, 32'h41737ec8};
test_label[2474] = '{32'h42001bd5};
test_output[2474] = '{32'h4260d538};
/*############ DEBUG ############
test_input[19792:19799] = '{32.027178426, -97.9242881748, 88.2354011282, 65.7566831416, 66.0058924035, -40.3392322725, 18.1137673336, 15.2184525474};
test_label[2474] = '{32.027178426};
test_output[2474] = '{56.2082227025};
############ END DEBUG ############*/
test_input[19800:19807] = '{32'hc1b7d09d, 32'h42554a14, 32'h42617323, 32'hc24de1fe, 32'hc292db27, 32'hc1c9617c, 32'hc2681a8d, 32'hc1fcb0d3};
test_label[2475] = '{32'hc1fcb0d3};
test_output[2475] = '{32'h42affdb2};
/*############ DEBUG ############
test_input[19800:19807] = '{-22.9768618605, 53.3223426442, 56.3624389551, -51.4706955041, -73.4280284558, -25.1725992568, -58.025930025, -31.5863408955};
test_label[2475] = '{-31.5863408955};
test_output[2475] = '{87.9955014794};
############ END DEBUG ############*/
test_input[19808:19815] = '{32'hc2a1e2d4, 32'hc2716d4e, 32'h429aae35, 32'h426807a1, 32'hc259a332, 32'hc2b06b1a, 32'hc292232d, 32'hc1fc1446};
test_label[2476] = '{32'h426807a1};
test_output[2476] = '{32'h419aa993};
/*############ DEBUG ############
test_input[19808:19815] = '{-80.9430238125, -60.3567445358, 77.340250493, 58.0074513421, -54.4093717388, -88.2091815192, -73.0687063553, -31.509899729};
test_label[2476] = '{58.0074513421};
test_output[2476] = '{19.3327991549};
############ END DEBUG ############*/
test_input[19816:19823] = '{32'h42632116, 32'hc2188f13, 32'h425056d4, 32'h4132920c, 32'h42857ade, 32'h411bcc5e, 32'hc1f1eeaf, 32'h41c49878};
test_label[2477] = '{32'hc1f1eeaf};
test_output[2477] = '{32'h42c1f690};
/*############ DEBUG ############
test_input[19816:19823] = '{56.7823113667, -38.1397213063, 52.0847940237, 11.1606556461, 66.7399763418, 9.73739416029, -30.2415440314, 24.5744477339};
test_label[2477] = '{-30.2415440314};
test_output[2477] = '{96.9815681671};
############ END DEBUG ############*/
test_input[19824:19831] = '{32'hc2967e71, 32'h42c62029, 32'h428e70f6, 32'hc15318d4, 32'hc28b404e, 32'h42204be4, 32'h428ce720, 32'h428cd467};
test_label[2478] = '{32'h428cd467};
test_output[2478] = '{32'h41e52f08};
/*############ DEBUG ############
test_input[19824:19831] = '{-75.2469589685, 99.0628139356, 71.220629092, -13.1935615446, -69.6255918967, 40.0741114357, 70.4514156812, 70.4148490886};
test_label[2478] = '{70.4148490886};
test_output[2478] = '{28.647964847};
############ END DEBUG ############*/
test_input[19832:19839] = '{32'hc2c2155b, 32'h429127bc, 32'h416ea517, 32'h40d0867a, 32'h42c4bd62, 32'h42c42170, 32'hc240d46c, 32'hc18ac771};
test_label[2479] = '{32'hc240d46c};
test_output[2479] = '{32'h43132137};
/*############ DEBUG ############
test_input[19832:19839] = '{-97.0417092759, 72.5776084647, 14.9153052453, 6.51641575766, 98.369887687, 98.0653084275, -48.2074425192, -17.347382657};
test_label[2479] = '{-48.2074425192};
test_output[2479] = '{147.129739275};
############ END DEBUG ############*/
test_input[19840:19847] = '{32'hc1f30ec1, 32'h4252138b, 32'h42b977d5, 32'hc2398002, 32'hc1a2c0a3, 32'hc223b1fa, 32'hc27bfc4f, 32'hc2683066};
test_label[2480] = '{32'hc2683066};
test_output[2480] = '{32'h4316c804};
/*############ DEBUG ############
test_input[19840:19847] = '{-30.3822033078, 52.5190867227, 92.7340432822, -46.3750074092, -20.3440615883, -40.9238064342, -62.9963950501, -58.0472651925};
test_label[2480] = '{-58.0472651925};
test_output[2480] = '{150.781308475};
############ END DEBUG ############*/
test_input[19848:19855] = '{32'hc25f2a91, 32'h42c06a17, 32'h419230e2, 32'h42c5f1f4, 32'hc18ffbc6, 32'h41dcdf8c, 32'h4040b07f, 32'hc287522b};
test_label[2481] = '{32'hc18ffbc6};
test_output[2481] = '{32'h42ea1028};
/*############ DEBUG ############
test_input[19848:19855] = '{-55.7915697328, 96.2072104908, 18.2738690897, 98.9725641578, -17.997937155, 27.609153798, 3.01077245117, -67.6604861287};
test_label[2481] = '{-17.997937155};
test_output[2481] = '{117.031552978};
############ END DEBUG ############*/
test_input[19856:19863] = '{32'h41131197, 32'h40fd3f98, 32'hc1a9dfee, 32'hc0baec0f, 32'hc1fdaf80, 32'hc22bc77c, 32'hc2b33a6e, 32'hc2a7b842};
test_label[2482] = '{32'hc1fdaf80};
test_output[2482] = '{32'h422497db};
/*############ DEBUG ############
test_input[19856:19863] = '{9.19179397785, 7.91401271248, -21.2343408908, -5.84131558264, -31.7106935244, -42.9448099265, -89.6141182818, -83.8598817999};
test_label[2482] = '{-31.7106935244};
test_output[2482] = '{41.1482963812};
############ END DEBUG ############*/
test_input[19864:19871] = '{32'h41788542, 32'hc2b15f1e, 32'h42994464, 32'hc1a09a7b, 32'h4264361d, 32'hc2af8f48, 32'h428e3ea1, 32'h42be64db};
test_label[2483] = '{32'hc2b15f1e};
test_output[2483] = '{32'h4337e1fc};
/*############ DEBUG ############
test_input[19864:19871] = '{15.5325339897, -88.6857766319, 76.6335743425, -20.0754290033, 57.0528443497, -87.7798461973, 71.1223183849, 95.1969824454};
test_label[2483] = '{-88.6857766319};
test_output[2483] = '{183.882759086};
############ END DEBUG ############*/
test_input[19872:19879] = '{32'h428180dd, 32'h424ba66c, 32'hc22fdd96, 32'hc2b6e5a7, 32'h4202c661, 32'hc1b32181, 32'hc26c9cd7, 32'hc0bce4e3};
test_label[2484] = '{32'hc26c9cd7};
test_output[2484] = '{32'h42f7cf49};
/*############ DEBUG ############
test_input[19872:19879] = '{64.7516872085, 50.9125225914, -43.966392736, -91.4485431728, 32.6937298638, -22.391358809, -59.1531623769, -5.90294028758};
test_label[2484] = '{-59.1531623769};
test_output[2484] = '{123.904850562};
############ END DEBUG ############*/
test_input[19880:19887] = '{32'h42bfae16, 32'hc2a98b4e, 32'h42334fcc, 32'h42271c4b, 32'hc2895a28, 32'h42805ad8, 32'h41af1ad4, 32'h4211dcdf};
test_label[2485] = '{32'h42271c4b};
test_output[2485] = '{32'h42583fe1};
/*############ DEBUG ############
test_input[19880:19887] = '{95.8400127293, -84.7720800657, 44.8279267164, 41.7776303467, -68.6760886918, 64.1774272224, 21.8881000177, 36.465693716};
test_label[2485] = '{41.7776303467};
test_output[2485] = '{54.0623823827};
############ END DEBUG ############*/
test_input[19888:19895] = '{32'h42741c2a, 32'hc028498d, 32'h4220406e, 32'h4291ff0c, 32'h4264cdd0, 32'h429ed140, 32'h424c9602, 32'hc257576d};
test_label[2486] = '{32'hc257576d};
test_output[2486] = '{32'h43053ee7};
/*############ DEBUG ############
test_input[19888:19895] = '{61.0275030409, -2.62948929634, 40.0629211968, 72.9981396307, 57.200987095, 79.4086922802, 51.146492271, -53.8353751049};
test_label[2486] = '{-53.8353751049};
test_output[2486] = '{133.245710161};
############ END DEBUG ############*/
test_input[19896:19903] = '{32'h41049977, 32'hc2bc1178, 32'hc0a6d0e8, 32'h42a5bd48, 32'hc2c7554d, 32'h41f0acfa, 32'h42a5fa3e, 32'h413da2d7};
test_label[2487] = '{32'hc2bc1178};
test_output[2487] = '{32'h4331a884};
/*############ DEBUG ############
test_input[19896:19903] = '{8.28746691115, -94.0341218619, -5.21300117464, 82.8696900727, -99.6666036971, 30.0844602865, 82.9887545742, 11.8522557963};
test_label[2487] = '{-94.0341218619};
test_output[2487] = '{177.658262365};
############ END DEBUG ############*/
test_input[19904:19911] = '{32'h42c2b149, 32'hbf6d1a32, 32'hc1fdb804, 32'hc1b2e4de, 32'h427a57ab, 32'h42842a68, 32'hc233eeed, 32'hc23a9c1b};
test_label[2488] = '{32'hc23a9c1b};
test_output[2488] = '{32'h430fffab};
/*############ DEBUG ############
test_input[19904:19911] = '{97.346261114, -0.926180957014, -31.7148516893, -22.3617511632, 62.58561243, 66.0828271856, -44.9833262004, -46.6524476704};
test_label[2488] = '{-46.6524476704};
test_output[2488] = '{143.998708784};
############ END DEBUG ############*/
test_input[19912:19919] = '{32'hc0d2b409, 32'hc22a8fc1, 32'hc2c672df, 32'hc24221d2, 32'h42a7af5b, 32'hc1f8c675, 32'hc269942b, 32'h41dbe346};
test_label[2489] = '{32'h41dbe346};
test_output[2489] = '{32'h42616d13};
/*############ DEBUG ############
test_input[19912:19919] = '{-6.58447711684, -42.6403846759, -99.2243610851, -48.5330286878, 83.8424896447, -31.0969024495, -58.3946939303, 27.4859736327};
test_label[2489] = '{27.4859736327};
test_output[2489] = '{56.3565160119};
############ END DEBUG ############*/
test_input[19920:19927] = '{32'hc1e74c60, 32'hc29d14d0, 32'h41a0828a, 32'hc197e197, 32'hc08d9969, 32'hc2b7a74c, 32'h4177f45f, 32'hbed9b464};
test_label[2490] = '{32'hc2b7a74c};
test_output[2490] = '{32'h42dfcd3a};
/*############ DEBUG ############
test_input[19920:19927] = '{-28.9122918622, -78.5406472561, 20.0637392795, -18.9851512919, -4.42497679495, -91.8267535273, 15.4971609142, -0.425204398387};
test_label[2490] = '{-91.8267535273};
test_output[2490] = '{111.900832629};
############ END DEBUG ############*/
test_input[19928:19935] = '{32'hc23701d7, 32'hc1d536ef, 32'h4294ec44, 32'h41c3fce9, 32'h427ee593, 32'h41813e28, 32'hc27430fe, 32'h428a9223};
test_label[2491] = '{32'hc1d536ef};
test_output[2491] = '{32'h42ca3ce5};
/*############ DEBUG ############
test_input[19928:19935] = '{-45.7517953093, -26.6518231466, 74.4614560193, 24.4984908393, 63.7241931527, 16.1553498189, -61.047842374, 69.2854249186};
test_label[2491] = '{-26.6518231466};
test_output[2491] = '{101.118935248};
############ END DEBUG ############*/
test_input[19936:19943] = '{32'hc296ce32, 32'hc26168c1, 32'hc113cc8b, 32'h41eee209, 32'hc226b0ae, 32'hc2c7f90f, 32'hc24f4b69, 32'h4226c2d7};
test_label[2492] = '{32'h41eee209};
test_output[2492] = '{32'h413d4753};
/*############ DEBUG ############
test_input[19936:19943] = '{-75.4027233798, -56.3522974094, -9.23743743636, 29.860369298, -41.6725381586, -99.9864407739, -51.8236435722, 41.6902749053};
test_label[2492] = '{29.860369298};
test_output[2492] = '{11.8299128908};
############ END DEBUG ############*/
test_input[19944:19951] = '{32'h41c0e7ad, 32'h422a6932, 32'h40e17c68, 32'hc2139a28, 32'h42043479, 32'hc2973bb9, 32'h41a79716, 32'h427f2b99};
test_label[2493] = '{32'h41a79716};
test_output[2493] = '{32'h422b600e};
/*############ DEBUG ############
test_input[19944:19951] = '{24.1131233067, 42.6027294837, 7.04643635254, -36.9005442716, 33.0512409536, -75.6166440555, 20.9487716388, 63.7925744727};
test_label[2493] = '{20.9487716388};
test_output[2493] = '{42.8438028345};
############ END DEBUG ############*/
test_input[19952:19959] = '{32'hc2c3283b, 32'hc201fef2, 32'h4266bd88, 32'h42040f91, 32'h414a219b, 32'h420a2c69, 32'h429cab3c, 32'hc2c7afc0};
test_label[2494] = '{32'hc201fef2};
test_output[2494] = '{32'h42ddaab5};
/*############ DEBUG ############
test_input[19952:19959] = '{-97.5785783759, -32.4989717039, 57.6850883439, 33.0152017556, 12.6332040885, 34.5433708007, 78.3344436275, -99.8432609422};
test_label[2494] = '{-32.4989717039};
test_output[2494] = '{110.833415332};
############ END DEBUG ############*/
test_input[19960:19967] = '{32'h4230dfa6, 32'hc119a8e5, 32'hc173ccc2, 32'h427f59f6, 32'hc1d30704, 32'h40cd8d1b, 32'hc1cafc1d, 32'h42063767};
test_label[2495] = '{32'h427f59f6};
test_output[2495] = '{32'h314f3d64};
/*############ DEBUG ############
test_input[19960:19967] = '{44.2184063841, -9.60373435627, -15.2374898445, 63.8378516632, -26.3784251516, 6.42347462086, -25.3731021034, 33.5541043223};
test_label[2495] = '{63.8378516632};
test_output[2495] = '{3.01573610983e-09};
############ END DEBUG ############*/
test_input[19968:19975] = '{32'h4281e04d, 32'h4289d4fa, 32'hc291385a, 32'hc1563580, 32'h4174c94c, 32'hc22d522f, 32'hc2b080de, 32'h42b51ec4};
test_label[2496] = '{32'hc2b080de};
test_output[2496] = '{32'h4332cfd1};
/*############ DEBUG ############
test_input[19968:19975] = '{64.9380893243, 68.9159675391, -72.6100609699, -13.3880615531, 15.2991444736, -43.3302587532, -88.2516901788, 90.5600858866};
test_label[2496] = '{-88.2516901788};
test_output[2496] = '{178.811776066};
############ END DEBUG ############*/
test_input[19976:19983] = '{32'h4287511d, 32'h423d25b0, 32'hc1a891a1, 32'h424744a7, 32'h42427063, 32'hc2a4780a, 32'h422cdfba, 32'hc29d6034};
test_label[2497] = '{32'h42427063};
test_output[2497] = '{32'h419863af};
/*############ DEBUG ############
test_input[19976:19983] = '{67.6584274306, 47.2868060403, -21.0711075679, 49.8170447587, 48.6097538288, -82.2344493777, 43.2184813725, -78.6878965305};
test_label[2497] = '{48.6097538288};
test_output[2497] = '{19.0486736264};
############ END DEBUG ############*/
test_input[19984:19991] = '{32'hc2c20d92, 32'hc2a1c25e, 32'h42c08ec5, 32'h42862431, 32'h421cbf21, 32'hc29c8229, 32'h42c1bd9a, 32'hc1b6a93f};
test_label[2498] = '{32'hc29c8229};
test_output[2498] = '{32'h432f90a8};
/*############ DEBUG ############
test_input[19984:19991] = '{-97.0265044898, -80.8796263764, 96.2788490876, 67.0706839551, 39.186648619, -78.2542179774, 96.870319206, -22.8326400464};
test_label[2498] = '{-78.2542179774};
test_output[2498] = '{175.565055974};
############ END DEBUG ############*/
test_input[19992:19999] = '{32'h429f212c, 32'h411a57c0, 32'hc2906f71, 32'hc0a89ff0, 32'h4220644d, 32'hc1fee460, 32'hc2a9ee1f, 32'h4281f3d4};
test_label[2499] = '{32'h4220644d};
test_output[2499] = '{32'h421dde0b};
/*############ DEBUG ############
test_input[19992:19999] = '{79.5647879713, 9.64642369667, -72.2176570989, -5.26952346504, 40.0979494875, -31.8615104253, -84.9650817012, 64.976229686};
test_label[2499] = '{40.0979494875};
test_output[2499] = '{39.4668389454};
############ END DEBUG ############*/
test_input[20000:20007] = '{32'hc2516151, 32'h41b64a6b, 32'hc2bcc21d, 32'hc22e2bcf, 32'h42829d46, 32'h41be132d, 32'h422a46cc, 32'h42839a67};
test_label[2500] = '{32'hc22e2bcf};
test_output[2500] = '{32'h42dba41f};
/*############ DEBUG ############
test_input[20000:20007] = '{-52.3450347636, 22.7863370805, -94.3791296992, -43.5427829422, 65.3071710226, 23.7593638506, 42.5691391998, 65.801566979};
test_label[2500] = '{-43.5427829422};
test_output[2500] = '{109.820546352};
############ END DEBUG ############*/
test_input[20008:20015] = '{32'hc14785c3, 32'h41bedad6, 32'hc22d8a71, 32'hc1c06e62, 32'h42b4b135, 32'h41d483c4, 32'h42154a52, 32'hc20c9a23};
test_label[2501] = '{32'h42154a52};
test_output[2501] = '{32'h42541818};
/*############ DEBUG ############
test_input[20008:20015] = '{-12.4701569257, 23.8568532143, -43.3851978435, -24.053898126, 90.3461100323, 26.5643387947, 37.3225798371, -35.1505230771};
test_label[2501] = '{37.3225798371};
test_output[2501] = '{53.0235301951};
############ END DEBUG ############*/
test_input[20016:20023] = '{32'h427e1563, 32'hc0cb840e, 32'h423664b3, 32'hc2ac901b, 32'hc1a4e9c3, 32'hc25f4be5, 32'hc1b881b9, 32'hc2a6e694};
test_label[2502] = '{32'h427e1563};
test_output[2502] = '{32'h328d5c3c};
/*############ DEBUG ############
test_input[20016:20023] = '{63.5208840434, -6.3598701311, 45.5983389647, -86.2814566588, -20.6141410416, -55.8241159814, -23.063341911, -83.4503510468};
test_label[2502] = '{63.5208840434};
test_output[2502] = '{1.64565036287e-08};
############ END DEBUG ############*/
test_input[20024:20031] = '{32'h41dc9daa, 32'h424aac92, 32'h41a9870c, 32'h4158719f, 32'h42a34390, 32'hc2b294f9, 32'hc1cc60d9, 32'hc2a63aff};
test_label[2503] = '{32'hc2a63aff};
test_output[2503] = '{32'h4324bf48};
/*############ DEBUG ############
test_input[20024:20031] = '{27.5769847315, 50.6685268673, 21.1909405795, 13.527739696, 81.6319567811, -89.2909628922, -25.5472886176, -83.1152296504};
test_label[2503] = '{-83.1152296504};
test_output[2503] = '{164.747186432};
############ END DEBUG ############*/
test_input[20032:20039] = '{32'h42aa803e, 32'h423efc29, 32'hc20795a3, 32'hc1d544dd, 32'h427da93c, 32'hc20f4856, 32'h42acbb4c, 32'h41cd3da2};
test_label[2504] = '{32'h42aa803e};
test_output[2504] = '{32'h3fb30e01};
/*############ DEBUG ############
test_input[20032:20039] = '{85.2504741248, 47.7462504823, -33.8961305615, -26.6586239463, 63.4152670414, -35.8206391876, 86.3658122693, 25.6550932945};
test_label[2504] = '{85.2504741248};
test_output[2504] = '{1.39886490689};
############ END DEBUG ############*/
test_input[20040:20047] = '{32'h429608b9, 32'hbfee6c13, 32'h4227d999, 32'h4289d477, 32'h42259a2b, 32'h3fa0a30d, 32'h42a67550, 32'hbfdf9dda};
test_label[2505] = '{32'h3fa0a30d};
test_output[2505] = '{32'h42a3f2e7};
/*############ DEBUG ############
test_input[20040:20047] = '{75.0170380182, -1.86267320206, 41.9624978603, 68.9149711653, 41.4005543368, 1.25497595608, 83.2291225946, -1.74700478983};
test_label[2505] = '{1.25497595608};
test_output[2505] = '{81.9744185633};
############ END DEBUG ############*/
test_input[20048:20055] = '{32'h42a7ced0, 32'hc2907a1f, 32'hc231b7ee, 32'h4238ed95, 32'hc2adff94, 32'h42a10922, 32'h42c27e98, 32'h400377db};
test_label[2506] = '{32'hc2907a1f};
test_output[2506] = '{32'h43297c5b};
/*############ DEBUG ############
test_input[20048:20055] = '{83.9039309704, -72.2385148438, -44.4296189576, 46.2320150822, -86.999177353, 80.5178385508, 97.2472528496, 2.05419032734};
test_label[2506] = '{-72.2385148438};
test_output[2506] = '{169.485769351};
############ END DEBUG ############*/
test_input[20056:20063] = '{32'h419e3964, 32'hc2074cad, 32'hc21c2b16, 32'hc231c476, 32'hc2613334, 32'hc2715cdb, 32'h406f55cc, 32'h42854c80};
test_label[2507] = '{32'h419e3964};
test_output[2507] = '{32'h423b7c4e};
/*############ DEBUG ############
test_input[20056:20063] = '{19.778021917, -33.8248804451, -39.0420752166, -44.4418571692, -56.3000017604, -60.3406779792, 3.73961154942, 66.6494139187};
test_label[2507] = '{19.778021917};
test_output[2507] = '{46.8713920017};
############ END DEBUG ############*/
test_input[20064:20071] = '{32'hc28f5c06, 32'hc1f25c75, 32'h418531bb, 32'h40c3917b, 32'hc232e996, 32'h4263eec1, 32'h42c25878, 32'h42628d11};
test_label[2508] = '{32'hc232e996};
test_output[2508] = '{32'h430de6a1};
/*############ DEBUG ############
test_input[20064:20071] = '{-71.6797361155, -30.2951456436, 16.6492815106, 6.11150890788, -44.7281102769, 56.9831576669, 97.1727893482, 56.6377616066};
test_label[2508] = '{-44.7281102769};
test_output[2508] = '{141.900899625};
############ END DEBUG ############*/
test_input[20072:20079] = '{32'hc2683477, 32'hc27c5815, 32'hc2bda404, 32'hc23ddccb, 32'hc2970b40, 32'hc1c672ee, 32'hbf9184ea, 32'h4234d4b7};
test_label[2509] = '{32'hc2bda404};
test_output[2509] = '{32'h430c0730};
/*############ DEBUG ############
test_input[20072:20079] = '{-58.0512361583, -63.0860172084, -94.8203422595, -47.4656162453, -75.5219732526, -24.8061186132, -1.13686870563, 45.2077296382};
test_label[2509] = '{-94.8203422595};
test_output[2509] = '{140.028071898};
############ END DEBUG ############*/
test_input[20080:20087] = '{32'h422d45d7, 32'hc203f28f, 32'hc2b6d059, 32'h4246bc14, 32'hc2b45a03, 32'hc2c312a3, 32'h41e36d3c, 32'hc2c07bb0};
test_label[2510] = '{32'hc2b45a03};
test_output[2510] = '{32'h430bdc77};
/*############ DEBUG ############
test_input[20080:20087] = '{43.3182031382, -32.986873546, -91.4069263531, 49.683671268, -90.175807845, -97.5364035359, 28.4283372037, -96.2415781991};
test_label[2510] = '{-90.175807845};
test_output[2510] = '{139.861197572};
############ END DEBUG ############*/
test_input[20088:20095] = '{32'hc2758603, 32'h42aefe1c, 32'h42abfb94, 32'hc291b76d, 32'h421bacff, 32'hc096c4dd, 32'h4296f794, 32'h42589cae};
test_label[2511] = '{32'h421bacff};
test_output[2511] = '{32'h42431c8e};
/*############ DEBUG ############
test_input[20088:20095] = '{-61.3808690017, 87.4963095616, 85.9913604636, -72.8582534964, 38.918939769, -4.71153113284, 75.4835528223, 54.1530065481};
test_label[2511] = '{38.918939769};
test_output[2511] = '{48.7778870176};
############ END DEBUG ############*/
test_input[20096:20103] = '{32'h424bc686, 32'h4287172c, 32'hc281a901, 32'h4213194e, 32'hc23acaf9, 32'h42c2fa91, 32'hc2a3fcbf, 32'hc22e29d6};
test_label[2512] = '{32'h424bc686};
test_output[2512] = '{32'h423a2e9c};
/*############ DEBUG ############
test_input[20096:20103] = '{50.9438695156, 67.5452550784, -64.8300875089, 36.7747120494, -46.6982149736, 97.4893852262, -81.9936482368, -43.5408566434};
test_label[2512] = '{50.9438695156};
test_output[2512] = '{46.5455157106};
############ END DEBUG ############*/
test_input[20104:20111] = '{32'hc2906f37, 32'h4287c977, 32'hc15156b0, 32'hc17e8d9d, 32'h428b540b, 32'hc232839b, 32'hc24b510f, 32'h41d3224f};
test_label[2513] = '{32'hc17e8d9d};
test_output[2513] = '{32'h42ab763a};
/*############ DEBUG ############
test_input[20104:20111] = '{-72.2172136848, 67.8934852261, -13.0836640806, -15.9095734818, 69.6641477886, -44.6285207501, -50.8291590489, 26.3917527921};
test_label[2513] = '{-15.9095734818};
test_output[2513] = '{85.7309131809};
############ END DEBUG ############*/
test_input[20112:20119] = '{32'hc2262b5d, 32'h42885b95, 32'h42865ccb, 32'h42ba9533, 32'h41158ab2, 32'h41509885, 32'hc28fd485, 32'hc2bc0a22};
test_label[2514] = '{32'h42885b95};
test_output[2514] = '{32'h41c8e676};
/*############ DEBUG ############
test_input[20112:20119] = '{-41.5423465564, 68.1788716645, 67.1812325357, 93.291401157, 9.34636077368, 13.0372357923, -71.9150787949, -94.0197885778};
test_label[2514] = '{68.1788716645};
test_output[2514] = '{25.1125294925};
############ END DEBUG ############*/
test_input[20120:20127] = '{32'h40a03ad7, 32'h427ecc2f, 32'h42c05fe2, 32'hc251d420, 32'h40ec92b3, 32'hc29325fd, 32'h41f4d3df, 32'hc2805c7f};
test_label[2515] = '{32'h42c05fe2};
test_output[2515] = '{32'h280c0000};
/*############ DEBUG ############
test_input[20120:20127] = '{5.00718258532, 63.6993974656, 96.187272645, -52.4571528481, 7.39290776145, -73.5741947272, 30.6034532771, -64.1806537991};
test_label[2515] = '{96.187272645};
test_output[2515] = '{7.77156117238e-15};
############ END DEBUG ############*/
test_input[20128:20135] = '{32'h4116c909, 32'hc201e799, 32'h425b0c4e, 32'h42af498f, 32'hc2ad03e7, 32'hc1cf48ec, 32'h422eaee7, 32'hc2a2564f};
test_label[2516] = '{32'hc1cf48ec};
test_output[2516] = '{32'h42e31bca};
/*############ DEBUG ############
test_input[20128:20135] = '{9.42408092621, -32.4761693608, 54.7620177313, 87.6436726576, -86.5076239043, -25.9106057816, 43.6708015082, -81.168575153};
test_label[2516] = '{-25.9106057816};
test_output[2516] = '{113.554278439};
############ END DEBUG ############*/
test_input[20136:20143] = '{32'hc24a0428, 32'h41f03525, 32'hc1ac3b62, 32'h427aefb8, 32'h423e30b3, 32'h41d5bd1a, 32'h41ce8ae0, 32'h41e872a8};
test_label[2517] = '{32'h41f03525};
test_output[2517] = '{32'h4202d525};
/*############ DEBUG ############
test_input[20136:20143] = '{-50.5040597507, 30.0259501691, -21.5289955927, 62.7341003834, 47.5475594473, 26.7173342546, 25.8178097551, 29.0559839763};
test_label[2517] = '{30.0259501691};
test_output[2517] = '{32.7081504681};
############ END DEBUG ############*/
test_input[20144:20151] = '{32'hc189293e, 32'h426687c6, 32'h42a3ce9a, 32'h4196685f, 32'h4202f0f1, 32'h421ab5c5, 32'hc1c44c6c, 32'hc19b6171};
test_label[2518] = '{32'h4196685f};
test_output[2518] = '{32'h427c6905};
/*############ DEBUG ############
test_input[20144:20151] = '{-17.145137848, 57.6325901262, 81.9035202504, 18.8009624353, 32.7352952607, 38.6775092015, -24.5373155533, -19.4225782134};
test_label[2518] = '{18.8009624353};
test_output[2518] = '{63.1025578151};
############ END DEBUG ############*/
test_input[20152:20159] = '{32'h41e61c8a, 32'hc0f56a6b, 32'hc283d75e, 32'h42c3318f, 32'hbe61ed8c, 32'h42bdcc42, 32'h41e12f1c, 32'h423a44e5};
test_label[2519] = '{32'h41e12f1c};
test_output[2519] = '{32'h428b0727};
/*############ DEBUG ############
test_input[20152:20159] = '{28.7639350099, -7.66924042251, -65.9206404895, 97.5967962941, -0.22063273875, 94.8989411834, 28.1480030707, 46.5672796877};
test_label[2519] = '{28.1480030707};
test_output[2519] = '{69.5139719919};
############ END DEBUG ############*/
test_input[20160:20167] = '{32'h42bc0c01, 32'h429d9d19, 32'h4246cff8, 32'h424edb1d, 32'h425095a8, 32'hc255fe0b, 32'h41b0de11, 32'hc292c5ea};
test_label[2520] = '{32'h429d9d19};
test_output[2520] = '{32'h4173773a};
/*############ DEBUG ############
test_input[20160:20167] = '{94.0234416061, 78.8068342068, 49.703095084, 51.7139761458, 52.1461481553, -53.4980885502, 22.1084302732, -73.3865544917};
test_label[2520] = '{78.8068342068};
test_output[2520] = '{15.2166076457};
############ END DEBUG ############*/
test_input[20168:20175] = '{32'h42bb03b2, 32'hc222e0f3, 32'h42b77b91, 32'h41a0bad7, 32'hc154b5a3, 32'h409312b1, 32'h42b36be0, 32'h42a96d8d};
test_label[2521] = '{32'h42b77b91};
test_output[2521] = '{32'h3ff8b082};
/*############ DEBUG ############
test_input[20168:20175] = '{93.5072202383, -40.7196773741, 91.7413379771, 20.0912304411, -13.2943452815, 4.59603179754, 89.710696003, 84.7139672466};
test_label[2521] = '{91.7413379771};
test_output[2521] = '{1.94288657131};
############ END DEBUG ############*/
test_input[20176:20183] = '{32'h41c787e9, 32'h42abda36, 32'hc2195c8d, 32'h42968eaa, 32'hc01ca76c, 32'h42bba187, 32'hc294a317, 32'hc2250f3e};
test_label[2522] = '{32'hc2250f3e};
test_output[2522] = '{32'h430714ac};
/*############ DEBUG ############
test_input[20176:20183] = '{24.9413620022, 85.9261927791, -38.3403824574, 75.2786438649, -2.44771858285, 93.8154827404, -74.3185320496, -41.2648863611};
test_label[2522] = '{-41.2648863611};
test_output[2522] = '{135.080743776};
############ END DEBUG ############*/
test_input[20184:20191] = '{32'hc2c0503d, 32'h41b5e537, 32'h42a45aa4, 32'hc1ab9162, 32'hc2b1dcee, 32'h423044df, 32'hc2803b9c, 32'h42966bb7};
test_label[2523] = '{32'h42966bb7};
test_output[2523] = '{32'h40def684};
/*############ DEBUG ############
test_input[20184:20191] = '{-96.156717544, 22.7369211594, 82.1770307664, -21.4459881922, -88.9315055089, 44.0672577731, -64.1164228661, 75.2103808362};
test_label[2523] = '{75.2103808362};
test_output[2523] = '{6.96759229214};
############ END DEBUG ############*/
test_input[20192:20199] = '{32'h414da4e3, 32'hc16a9809, 32'h42a5ef89, 32'h41e3eec3, 32'hc2be3c21, 32'hc1998a7a, 32'h41dae0b7, 32'h41bd6f48};
test_label[2524] = '{32'h41dae0b7};
test_output[2524] = '{32'h425e6eb6};
/*############ DEBUG ############
test_input[20192:20199] = '{12.8527554503, -14.6621183425, 82.9678398535, 28.4915827876, -95.1174399098, -19.192615636, 27.3597238014, 23.6793365003};
test_label[2524] = '{27.3597238014};
test_output[2524] = '{55.6081160521};
############ END DEBUG ############*/
test_input[20200:20207] = '{32'hc26ac36d, 32'h429bcc87, 32'hc20b6902, 32'h410e0e0c, 32'h423c046b, 32'hc29b1e58, 32'h425cfa7b, 32'h429cacb6};
test_label[2525] = '{32'hc29b1e58};
test_output[2525] = '{32'h431c6503};
/*############ DEBUG ############
test_input[20200:20207] = '{-58.6908443173, 77.8994661719, -34.852547359, 8.87842895752, 47.0043147199, -77.5592660957, 55.2446087136, 78.3373234821};
test_label[2525] = '{-77.5592660957};
test_output[2525] = '{156.394583955};
############ END DEBUG ############*/
test_input[20208:20215] = '{32'hc1465063, 32'h427b7fb7, 32'hc2bd2262, 32'h40d33d66, 32'h42608355, 32'hc295c8a1, 32'hc2a43eed, 32'h42c61389};
test_label[2526] = '{32'h42c61389};
test_output[2526] = '{32'h25800000};
/*############ DEBUG ############
test_input[20208:20215] = '{-12.3946257366, 62.8747228807, -94.5671546272, 6.60124479392, 56.1282532943, -74.8918501618, -82.1229051052, 99.0381543578};
test_label[2526] = '{99.0381543578};
test_output[2526] = '{2.22044604925e-16};
############ END DEBUG ############*/
test_input[20216:20223] = '{32'hc19aaa2c, 32'hc227ac90, 32'hc2c37547, 32'hc2bf44ea, 32'h41afc9b7, 32'h4286a71d, 32'hc16b4fd8, 32'h4257a75c};
test_label[2527] = '{32'h4257a75c};
test_output[2527] = '{32'h41569b79};
/*############ DEBUG ############
test_input[20216:20223] = '{-19.3330912887, -41.9185193, -97.7290538642, -95.6345971694, 21.9734942313, 67.3263915021, -14.70699314, 53.9134356264};
test_label[2527] = '{53.9134356264};
test_output[2527] = '{13.4129573713};
############ END DEBUG ############*/
test_input[20224:20231] = '{32'hc2bd7d61, 32'hc2870a93, 32'hc1bc818c, 32'hc2830f13, 32'hc0be478d, 32'h41f63368, 32'hc0d2fac7, 32'hc2278f95};
test_label[2528] = '{32'hc2278f95};
test_output[2528] = '{32'h429154a4};
/*############ DEBUG ############
test_input[20224:20231] = '{-94.7448769667, -67.5206535845, -23.5632557429, -65.5294421578, -5.94623405694, 30.7751007453, -6.59311245754, -41.8902166047};
test_label[2528] = '{-41.8902166047};
test_output[2528] = '{72.66531735};
############ END DEBUG ############*/
test_input[20232:20239] = '{32'hc2250f8b, 32'hc2872278, 32'h419de572, 32'h420fbc42, 32'h412dc155, 32'hc2bcf8c0, 32'h42a6eea6, 32'h3f84dfc2};
test_label[2529] = '{32'h420fbc42};
test_output[2529] = '{32'h423e210b};
/*############ DEBUG ############
test_input[20232:20239] = '{-41.2651801359, -67.567321516, 19.7370331712, 35.9338448097, 10.859700143, -94.485841789, 83.46611345, 1.03807853017};
test_label[2529] = '{35.9338448097};
test_output[2529] = '{47.5322686403};
############ END DEBUG ############*/
test_input[20240:20247] = '{32'h41511d51, 32'h42c3f08a, 32'h41b809de, 32'h4186b90a, 32'h42815fd2, 32'h42c2b8fc, 32'hc20173f7, 32'h42a6568e};
test_label[2530] = '{32'h42815fd2};
test_output[2530] = '{32'h4206de5a};
/*############ DEBUG ############
test_input[20240:20247] = '{13.0696576441, 97.9698011544, 23.00481771, 16.8403504616, 64.6871458022, 97.3612998981, -32.3632470377, 83.1690483229};
test_label[2530] = '{64.6871458022};
test_output[2530] = '{33.7171394383};
############ END DEBUG ############*/
test_input[20248:20255] = '{32'h423de2e9, 32'hc28a3d8d, 32'hc2ba042e, 32'hc241ba95, 32'hc28b5905, 32'h42bb55d3, 32'h428755f8, 32'hc2639e7e};
test_label[2531] = '{32'hc2ba042e};
test_output[2531] = '{32'h433aad00};
/*############ DEBUG ############
test_input[20248:20255] = '{47.4715934855, -69.1202156866, -93.0081627005, -48.4322101821, -69.6738657206, 93.6676261329, 67.6679095446, -56.9047771993};
test_label[2531] = '{-93.0081627005};
test_output[2531] = '{186.675788833};
############ END DEBUG ############*/
test_input[20256:20263] = '{32'hc296d1cb, 32'h41eaaf49, 32'h42521541, 32'h4086d428, 32'h419dc7f8, 32'h41b358a1, 32'hc1e42071, 32'hc1d3197e};
test_label[2532] = '{32'h41eaaf49};
test_output[2532] = '{32'h41b97b39};
/*############ DEBUG ############
test_input[20256:20263] = '{-75.4097494764, 29.3355883486, 52.520755852, 4.21339793044, 19.7226417945, 22.4182767797, -28.5158396022, -26.3874477911};
test_label[2532] = '{29.3355883486};
test_output[2532] = '{23.1851675035};
############ END DEBUG ############*/
test_input[20264:20271] = '{32'hc2aa491b, 32'h428d19bd, 32'h42af28fd, 32'h423a6b25, 32'hc2c0db96, 32'h42b1e0c8, 32'h41c85fe0, 32'h4299b4a2};
test_label[2533] = '{32'h423a6b25};
test_output[2533] = '{32'h422a4095};
/*############ DEBUG ############
test_input[20264:20271] = '{-85.1427830475, 70.5502701425, 87.580054392, 46.6046327628, -96.4288822975, 88.9390275516, 25.0468144642, 76.852801019};
test_label[2533] = '{46.6046327628};
test_output[2533] = '{42.5630671153};
############ END DEBUG ############*/
test_input[20272:20279] = '{32'hc2085635, 32'h4164c8c7, 32'h41a02515, 32'hc243aae0, 32'h416006c1, 32'hc20277bd, 32'h427d5831, 32'hc2908620};
test_label[2534] = '{32'h427d5831};
test_output[2534] = '{32'h80000000};
/*############ DEBUG ############
test_input[20272:20279] = '{-34.0841863446, 14.299018227, 20.0181058919, -48.9168698694, 14.0016491602, -32.6169323224, 63.3361260252, -72.2619609834};
test_label[2534] = '{63.3361260252};
test_output[2534] = '{-0.0};
############ END DEBUG ############*/
test_input[20280:20287] = '{32'h42b9465b, 32'hc2c72c1a, 32'hc16ee097, 32'hc2a5caf4, 32'hc0308858, 32'hc168d591, 32'hc2467e42, 32'hc208d273};
test_label[2535] = '{32'hc2a5caf4};
test_output[2535] = '{32'h432f88a8};
/*############ DEBUG ############
test_input[20280:20287] = '{92.637414891, -99.5861381387, -14.9298319129, -82.8963927898, -2.75832172001, -14.5521406889, -49.6232974394, -34.2055180792};
test_label[2535] = '{-82.8963927898};
test_output[2535] = '{175.533807681};
############ END DEBUG ############*/
test_input[20288:20295] = '{32'hc25aaa05, 32'hc2a595e2, 32'hc24bb46b, 32'hc210b9a8, 32'hc197f755, 32'hc219964a, 32'hc1c225b6, 32'hc1cd8a8c};
test_label[2536] = '{32'hc219964a};
test_output[2536] = '{32'h419b423e};
/*############ DEBUG ############
test_input[20288:20295] = '{-54.6660359047, -82.792736445, -50.9261890719, -36.1813041062, -18.9957679706, -38.3967683176, -24.2684138478, -25.6926490253};
test_label[2536] = '{-38.3967683176};
test_output[2536] = '{19.4073449915};
############ END DEBUG ############*/
test_input[20296:20303] = '{32'hc2a52f95, 32'hc2353fbf, 32'hc273bee9, 32'h428fb13d, 32'h40cba763, 32'hc2b82b81, 32'hc2b82dd4, 32'h42bbde90};
test_label[2537] = '{32'hc2353fbf};
test_output[2537] = '{32'h430b3f38};
/*############ DEBUG ############
test_input[20296:20303] = '{-82.5929352881, -45.3122504532, -60.9364343327, 71.8461686683, 6.36418295018, -92.0849683755, -92.0895101892, 93.9346906958};
test_label[2537] = '{-45.3122504532};
test_output[2537] = '{139.246941149};
############ END DEBUG ############*/
test_input[20304:20311] = '{32'hc2ba285d, 32'h42912410, 32'hc12a24e3, 32'hc26dd6b3, 32'hc07daa14, 32'hc2741a5b, 32'h417db784, 32'h4290c8bd};
test_label[2538] = '{32'hc2741a5b};
test_output[2538] = '{32'h43063440};
/*############ DEBUG ############
test_input[20304:20311] = '{-93.0788356807, 72.5704346104, -10.6340053092, -59.4596667627, -3.96350563038, -61.0257359578, 15.8573039785, 72.3920654906};
test_label[2538] = '{-61.0257359578};
test_output[2538] = '{134.204104871};
############ END DEBUG ############*/
test_input[20312:20319] = '{32'hc20ac129, 32'hc28322ea, 32'h412b9ba3, 32'h427ff130, 32'hc221a00e, 32'hc28fc624, 32'h423b4b9d, 32'h4214abaa};
test_label[2539] = '{32'h427ff130};
test_output[2539] = '{32'h33174599};
/*############ DEBUG ############
test_input[20312:20319] = '{-34.6886316144, -65.5681944302, 10.725497027, 63.9855362943, -40.4063051323, -71.8869924485, 46.8238411176, 37.1676404298};
test_label[2539] = '{63.9855362943};
test_output[2539] = '{3.52207244022e-08};
############ END DEBUG ############*/
test_input[20320:20327] = '{32'h421f3deb, 32'h42651d82, 32'hc164a009, 32'hc28871c4, 32'h41cfb53e, 32'hc17d52c8, 32'hc2c0bbc4, 32'h4243625f};
test_label[2540] = '{32'h41cfb53e};
test_output[2540] = '{32'h41fa8638};
/*############ DEBUG ############
test_input[20320:20327] = '{39.8104662199, 57.278816613, -14.2890713722, -68.2221995649, 25.9634979876, -15.8327100014, -96.3667275089, 48.8460641557};
test_label[2540] = '{25.9634979876};
test_output[2540] = '{31.3155362493};
############ END DEBUG ############*/
test_input[20328:20335] = '{32'hc2c5a790, 32'h427975e7, 32'h42336f21, 32'hc2227f4c, 32'h42b2f347, 32'h42953953, 32'h41a9cf6f, 32'hc094c3b2};
test_label[2541] = '{32'h42953953};
test_output[2541] = '{32'h416dcfa1};
/*############ DEBUG ############
test_input[20328:20335] = '{-98.827267511, 62.3651392514, 44.8585234218, -40.6243124291, 89.4751503996, 74.6119601074, 21.2262859791, -4.64888863221};
test_label[2541] = '{74.6119601074};
test_output[2541] = '{14.8631906429};
############ END DEBUG ############*/
test_input[20336:20343] = '{32'h424eb413, 32'hc2b524d9, 32'hc18cb55a, 32'h4249e61b, 32'h3ec4ba4b, 32'h41a17b55, 32'hc229f2ad, 32'hc2bdf79a};
test_label[2542] = '{32'h4249e61b};
test_output[2542] = '{32'h3fbb6991};
/*############ DEBUG ############
test_input[20336:20343] = '{51.6758530788, -90.5719714135, -17.5885508795, 50.4747125808, 0.384233794125, 20.1852213987, -42.486987108, -94.98359411};
test_label[2542] = '{50.4747125808};
test_output[2542] = '{1.46415908399};
############ END DEBUG ############*/
test_input[20344:20351] = '{32'h429ef1fa, 32'h3fbf5701, 32'hc2686d4b, 32'h427bbf62, 32'h4289b292, 32'h42737495, 32'hc2bb9d04, 32'hc2b301d5};
test_label[2543] = '{32'hc2bb9d04};
test_output[2543] = '{32'h432d4781};
/*############ DEBUG ############
test_input[20344:20351] = '{79.4726103256, 1.49484263212, -58.106732054, 62.9368985418, 68.8487671553, 60.8638480796, -93.8066703579, -89.5035743892};
test_label[2543] = '{-93.8066703579};
test_output[2543] = '{173.279305086};
############ END DEBUG ############*/
test_input[20352:20359] = '{32'h400da7c9, 32'hc2241ae4, 32'hc2c64a09, 32'h426891a5, 32'hc1032442, 32'h429a9122, 32'h428cf744, 32'hc280611a};
test_label[2544] = '{32'h426891a5};
test_output[2544] = '{32'h41992388};
/*############ DEBUG ############
test_input[20352:20359] = '{2.21336576079, -41.0262620278, -99.1445975186, 58.1422296427, -8.19635159979, 77.2834654903, 70.4829421785, -64.1896510497};
test_label[2544] = '{58.1422296427};
test_output[2544] = '{19.1423484259};
############ END DEBUG ############*/
test_input[20360:20367] = '{32'hc29e5401, 32'hc2a85d73, 32'h422e9f47, 32'h42869529, 32'hc28f429b, 32'h42bbc001, 32'h429a1066, 32'hc244fb1b};
test_label[2545] = '{32'hc28f429b};
test_output[2545] = '{32'h4325814e};
/*############ DEBUG ############
test_input[20360:20367] = '{-79.1640678293, -84.1825180628, 43.6555444941, 67.2913284346, -71.6300872707, 93.8750068243, 77.0320317063, -49.2452217525};
test_label[2545] = '{-71.6300872707};
test_output[2545] = '{165.505094143};
############ END DEBUG ############*/
test_input[20368:20375] = '{32'hc27911df, 32'h41462c47, 32'hbfdd01be, 32'h420cf551, 32'hc2bfa3fc, 32'hc283c70e, 32'hc2b4ced1, 32'hc2a2b5e0};
test_label[2546] = '{32'h41462c47};
test_output[2546] = '{32'h41b6d47f};
/*############ DEBUG ############
test_input[20368:20375] = '{-62.2674529593, 12.3858095153, -1.72661571664, 35.2395677594, -95.820281094, -65.8887816133, -90.4039415224, -81.3552230218};
test_label[2546] = '{12.3858095153};
test_output[2546] = '{22.8537582442};
############ END DEBUG ############*/
test_input[20376:20383] = '{32'hc2c0c85a, 32'h4280a717, 32'hc1858bae, 32'h41c0ea4c, 32'h4216e94c, 32'h423f46c0, 32'hc0d4c5d6, 32'hc1c2c3b7};
test_label[2547] = '{32'hc1c2c3b7};
test_output[2547] = '{32'h42b15805};
/*############ DEBUG ############
test_input[20376:20383] = '{-96.3913088421, 64.3263509956, -16.6932039256, 24.1144024874, 37.7278293351, 47.8190936913, -6.6491497756, -24.3455640461};
test_label[2547] = '{-24.3455640461};
test_output[2547] = '{88.6719151095};
############ END DEBUG ############*/
test_input[20384:20391] = '{32'h425c7ee4, 32'h420fcdbf, 32'h42231723, 32'h42bf34bf, 32'h42849b19, 32'hc281f856, 32'h4226324b, 32'hc2a5e97d};
test_label[2548] = '{32'hc2a5e97d};
test_output[2548] = '{32'h43328f1e};
/*############ DEBUG ############
test_input[20384:20391] = '{55.1239155054, 35.9509243792, 40.7725930577, 95.6030160779, 66.3029278976, -64.9850343977, 41.5491139301, -82.9560298062};
test_label[2548] = '{-82.9560298062};
test_output[2548] = '{178.559045884};
############ END DEBUG ############*/
test_input[20392:20399] = '{32'hc2b219a6, 32'h416b200e, 32'hc256dabf, 32'hc282ef65, 32'hc1f54aa2, 32'hc12ec380, 32'h426cc1d0, 32'hc289ede8};
test_label[2549] = '{32'hc289ede8};
test_output[2549] = '{32'h43002768};
/*############ DEBUG ############
test_input[20392:20399] = '{-89.0500951752, 14.6953261603, -53.713617581, -65.4675658571, -30.6614414548, -10.9227292816, 59.18926963, -68.9646622792};
test_label[2549] = '{-68.9646622792};
test_output[2549] = '{128.153931909};
############ END DEBUG ############*/
test_input[20400:20407] = '{32'h42313068, 32'h42c0a6c3, 32'hc1cfba4a, 32'hc29a85d5, 32'hc2a44cb2, 32'h41e7f6eb, 32'h429739a5, 32'hc2b6bd8c};
test_label[2550] = '{32'h42c0a6c3};
test_output[2550] = '{32'h308ad704};
/*############ DEBUG ############
test_input[20400:20407] = '{44.297271938, 96.3257097216, -25.9659619568, -77.2613894658, -82.1497952997, 28.9955649834, 75.6125855423, -91.3702105831};
test_label[2550] = '{96.3257097216};
test_output[2550] = '{1.01019326288e-09};
############ END DEBUG ############*/
test_input[20408:20415] = '{32'h4294627d, 32'h41880028, 32'hc2c6c8a2, 32'hc252be33, 32'hc281dca1, 32'h4216bae3, 32'hc20b83ff, 32'hc294f15c};
test_label[2551] = '{32'h4216bae3};
test_output[2551] = '{32'h42120a17};
/*############ DEBUG ############
test_input[20408:20415] = '{74.1923587121, 17.0000771539, -99.3918591113, -52.6857431849, -64.9309143429, 37.6825053831, -34.8789009061, -74.4714034952};
test_label[2551] = '{37.6825053831};
test_output[2551] = '{36.509853329};
############ END DEBUG ############*/
test_input[20416:20423] = '{32'hc23a9de1, 32'hc19b8e5b, 32'h41c3aa2a, 32'hc221607b, 32'h42609a6e, 32'h429b8f99, 32'h425f7668, 32'hc11da7e1};
test_label[2552] = '{32'hc23a9de1};
test_output[2552] = '{32'h42f8de8a};
/*############ DEBUG ############
test_input[20416:20423] = '{-46.6541787335, -19.4445096846, 24.4580883071, -40.3442182701, 56.1508088382, 77.7804661243, 55.865632149, -9.85348636831};
test_label[2552] = '{-46.6541787335};
test_output[2552] = '{124.434644859};
############ END DEBUG ############*/
test_input[20424:20431] = '{32'h42b4e5d0, 32'hc201ed92, 32'h427f0e7b, 32'hc245cf91, 32'hc253452d, 32'h422a3cb4, 32'h4266553b, 32'h42a9680a};
test_label[2553] = '{32'hc253452d};
test_output[2553] = '{32'h430f4504};
/*############ DEBUG ############
test_input[20424:20431] = '{90.4488513053, -32.4820008988, 63.7641410382, -49.4527025858, -52.8175558436, 42.5592819801, 57.5832345648, 84.7032014855};
test_label[2553] = '{-52.8175558436};
test_output[2553] = '{143.269598707};
############ END DEBUG ############*/
test_input[20432:20439] = '{32'hc2a6629a, 32'h427a8b78, 32'hc14317de, 32'hc178e9a7, 32'h41897e79, 32'hbd080438, 32'h4132017c, 32'h41f944a9};
test_label[2554] = '{32'hc178e9a7};
test_output[2554] = '{32'h429c62f1};
/*############ DEBUG ############
test_input[20432:20439] = '{-83.1925789121, 62.6361984577, -12.1933268901, -15.5570440402, 17.1867548788, -0.0332071497092, 11.1253624383, 31.1585261498};
test_label[2554] = '{-15.5570440402};
test_output[2554] = '{78.1932424979};
############ END DEBUG ############*/
test_input[20440:20447] = '{32'hc241ee84, 32'hc295580e, 32'h423118ba, 32'h4159c749, 32'h4096145c, 32'hc29399ae, 32'hc2c78306, 32'h428b8bdd};
test_label[2555] = '{32'h4096145c};
test_output[2555] = '{32'h42822a97};
/*############ DEBUG ############
test_input[20440:20447] = '{-48.4829250513, -74.671979238, 44.2741487548, 13.6111538624, 4.68998506419, -73.8001544725, -99.755904474, 69.7731671968};
test_label[2555] = '{4.68998506419};
test_output[2555] = '{65.0831821326};
############ END DEBUG ############*/
test_input[20448:20455] = '{32'hc18e4c6b, 32'h42063a04, 32'hc26c825b, 32'hc282e498, 32'hc152d0a8, 32'hc29cc1d3, 32'h41ee5534, 32'h42811ae6};
test_label[2556] = '{32'hc26c825b};
test_output[2556] = '{32'h42f75c13};
/*############ DEBUG ############
test_input[20448:20455] = '{-17.7873142499, 33.5566566328, -59.1272995412, -65.4464740159, -13.1759417094, -78.3785639798, 29.7916024652, 64.5525360331};
test_label[2556] = '{-59.1272995412};
test_output[2556] = '{123.679835574};
############ END DEBUG ############*/
test_input[20456:20463] = '{32'hc21106e8, 32'hc1e7fda0, 32'hc286e9cb, 32'hc1bb5671, 32'hc2707b9d, 32'hc28d7084, 32'hbfe81bb5, 32'h40a828bc};
test_label[2557] = '{32'hc2707b9d};
test_output[2557] = '{32'h4282c0ca};
/*############ DEBUG ############
test_input[20456:20463] = '{-36.2567442238, -28.9988398147, -67.4566272508, -23.4172081476, -60.1207145644, -70.7197557236, -1.81334559722, 5.25497242394};
test_label[2557] = '{-60.1207145644};
test_output[2557] = '{65.3765382903};
############ END DEBUG ############*/
test_input[20464:20471] = '{32'h424b8ce9, 32'hc0558c4c, 32'h42b44332, 32'hc29a1fbb, 32'hc11dc1a1, 32'hc2551aec, 32'h4128c8f7, 32'hc1a7e074};
test_label[2558] = '{32'hc11dc1a1};
test_output[2558] = '{32'h42c7fb66};
/*############ DEBUG ############
test_input[20464:20471] = '{50.8876092667, -3.33668815191, 90.1312420633, -77.0619718898, -9.85977276968, -53.2762927701, 10.5490633288, -20.9845953847};
test_label[2558] = '{-9.85977276968};
test_output[2558] = '{99.991014833};
############ END DEBUG ############*/
test_input[20472:20479] = '{32'hc28b7216, 32'h4248732d, 32'h42a5a89f, 32'h4151b5be, 32'hc28545d6, 32'hc290251d, 32'hc274fd09, 32'hc29dd678};
test_label[2559] = '{32'hc28b7216};
test_output[2559] = '{32'h43188d5b};
/*############ DEBUG ############
test_input[20472:20479] = '{-69.7228255411, 50.1124781505, 82.8293367289, 13.1068710526, -66.6363972362, -72.0724852006, -61.2471041062, -78.9188852387};
test_label[2559] = '{-69.7228255411};
test_output[2559] = '{152.55216227};
############ END DEBUG ############*/
test_input[20480:20487] = '{32'hc26b9be0, 32'h4184ad11, 32'hc20d9b29, 32'h420c29ab, 32'h428f0c24, 32'h42b5fca5, 32'hc254dbc0, 32'h41dc3f40};
test_label[2560] = '{32'h428f0c24};
test_output[2560] = '{32'h419bc205};
/*############ DEBUG ############
test_input[20480:20487] = '{-58.9022205641, 16.5845057827, -35.401522257, 35.0406927826, 71.5237092226, 90.993445765, -53.2146003041, 27.5308843776};
test_label[2560] = '{71.5237092226};
test_output[2560] = '{19.469736546};
############ END DEBUG ############*/
test_input[20488:20495] = '{32'h424be9a3, 32'hc1fcd834, 32'h428efac4, 32'hc0e06be0, 32'hc27bd358, 32'hc296028e, 32'hc20d2476, 32'hc2433e3e};
test_label[2561] = '{32'hc2433e3e};
test_output[2561] = '{32'h42f099e3};
/*############ DEBUG ############
test_input[20488:20495] = '{50.9781619707, -31.6055686781, 71.4897743342, -7.01316819926, -62.9563892464, -75.004993393, -35.2856081896, -48.8107843463};
test_label[2561] = '{-48.8107843463};
test_output[2561] = '{120.300558682};
############ END DEBUG ############*/
test_input[20496:20503] = '{32'h42a2708a, 32'h40f17e53, 32'hc2ae878f, 32'hc29bfd66, 32'hc2501ad4, 32'hc2496e37, 32'h428fc253, 32'hc244703f};
test_label[2562] = '{32'hc2496e37};
test_output[2562] = '{32'h430393d9};
/*############ DEBUG ############
test_input[20496:20503] = '{81.2198054544, 7.54667055035, -87.2647637827, -77.9949212411, -52.0261989653, -50.3576312375, 71.8795387092, -49.109614047};
test_label[2562] = '{-50.3576312375};
test_output[2562] = '{131.577524504};
############ END DEBUG ############*/
test_input[20504:20511] = '{32'hc2c2e0bf, 32'hc2a8dd67, 32'hc27fb518, 32'h41af347c, 32'h42ac701a, 32'h4170684e, 32'h41b72118, 32'hc16b07f9};
test_label[2563] = '{32'h41b72118};
test_output[2563] = '{32'h427d4fa8};
/*############ DEBUG ############
test_input[20504:20511] = '{-97.4389548241, -84.43242853, -63.9268481999, 21.9006262931, 86.2189469061, 15.0254652106, 22.8911587996, -14.6894466743};
test_label[2563] = '{22.8911587996};
test_output[2563] = '{63.3277881065};
############ END DEBUG ############*/
test_input[20512:20519] = '{32'hc28d80b8, 32'h4262c5aa, 32'h42a9230d, 32'hc2ade081, 32'hc1ac7c0b, 32'hbffc3eff, 32'h428ca428, 32'h42670a8b};
test_label[2564] = '{32'hc2ade081};
test_output[2564] = '{32'h432b81c7};
/*############ DEBUG ############
test_input[20512:20519] = '{-70.7514061181, 56.6930301847, 84.5684611542, -86.9384861636, -21.5605684974, -1.97067248185, 70.3206201176, 57.760295812};
test_label[2564] = '{-86.9384861636};
test_output[2564] = '{171.506947967};
############ END DEBUG ############*/
test_input[20520:20527] = '{32'h42a97496, 32'h42656451, 32'h41da0675, 32'h42ba49e0, 32'hc2992a56, 32'h4288b579, 32'hc0eee461, 32'hc23faf6c};
test_label[2565] = '{32'hc0eee461};
test_output[2565] = '{32'h42c93843};
/*############ DEBUG ############
test_input[20520:20527] = '{84.7277060852, 57.3479663518, 27.2531527358, 93.1442902041, -76.5826846847, 68.3544364573, -7.46537815977, -47.9213099471};
test_label[2565] = '{-7.46537815977};
test_output[2565] = '{100.609889508};
############ END DEBUG ############*/
test_input[20528:20535] = '{32'hc28ceb1f, 32'h41da3019, 32'h424371ac, 32'hc293e4d0, 32'h42c3621c, 32'hc1b2cf58, 32'h401833ff, 32'h42ab37f2};
test_label[2566] = '{32'h401833ff};
test_output[2566] = '{32'h42bea07d};
/*############ DEBUG ############
test_input[20528:20535] = '{-70.4592218894, 27.2734846399, 48.861008938, -73.9468999074, 97.6916204801, -22.3512415641, 2.37817356757, 85.6092716766};
test_label[2566] = '{2.37817356757};
test_output[2566] = '{95.313452571};
############ END DEBUG ############*/
test_input[20536:20543] = '{32'hc1fc1ea5, 32'h4296cd5c, 32'h42af4859, 32'hc2c5d5d9, 32'hc27db856, 32'hc231ac90, 32'hc2c7bab9, 32'h41c331e2};
test_label[2567] = '{32'h41c331e2};
test_output[2567] = '{32'h427cf7c2};
/*############ DEBUG ############
test_input[20536:20543] = '{-31.514963149, 75.401092148, 87.6413021608, -98.9176743106, -63.430015651, -44.4185176278, -99.8646902172, 24.399357127};
test_label[2567] = '{24.399357127};
test_output[2567] = '{63.2419498661};
############ END DEBUG ############*/
test_input[20544:20551] = '{32'hc09dda42, 32'hc20d18cb, 32'hc1896364, 32'h42c4c821, 32'h413015bf, 32'hc191a64a, 32'h42979a0b, 32'h42c0bbdc};
test_label[2568] = '{32'h42979a0b};
test_output[2568] = '{32'h41b5b67f};
/*############ DEBUG ############
test_input[20544:20551] = '{-4.93289272432, -35.2742137804, -17.173531158, 98.3908735399, 11.00530906, -18.2061953399, 75.8008656031, 96.3669162925};
test_label[2568] = '{75.8008656031};
test_output[2568] = '{22.7141101218};
############ END DEBUG ############*/
test_input[20552:20559] = '{32'hc29aa261, 32'h41e6e0c4, 32'hc2a49b0e, 32'h42138ee4, 32'h42080901, 32'hc2a05241, 32'h4132ec01, 32'h422b8cab};
test_label[2569] = '{32'h41e6e0c4};
test_output[2569] = '{32'h41607be2};
/*############ DEBUG ############
test_input[20552:20559] = '{-77.3171473508, 28.8597483797, -82.3028432857, 36.8895400696, 34.0087934481, -80.1606550097, 11.1826176995, 42.8873723622};
test_label[2569] = '{28.8597483797};
test_output[2569] = '{14.0302448271};
############ END DEBUG ############*/
test_input[20560:20567] = '{32'hc2370824, 32'hc267fdd5, 32'h423cf73c, 32'hc23f2891, 32'h42110862, 32'h42ba47bc, 32'hc1adc0a1, 32'hc2c50493};
test_label[2570] = '{32'hc1adc0a1};
test_output[2570] = '{32'h42e5b7e4};
/*############ DEBUG ############
test_input[20560:20567] = '{-45.7579484199, -57.9978827715, 47.2414395615, -47.7896171558, 36.2581864941, 93.1401054015, -21.7190564395, -98.5089340704};
test_label[2570] = '{-21.7190564395};
test_output[2570] = '{114.859161841};
############ END DEBUG ############*/
test_input[20568:20575] = '{32'hc1c445a3, 32'h4203f655, 32'h42891c6a, 32'h428a569e, 32'h4215590a, 32'h425148b6, 32'h4285efa1, 32'hbf52e85d};
test_label[2571] = '{32'h428a569e};
test_output[2571] = '{32'h3f008377};
/*############ DEBUG ############
test_input[20568:20575] = '{-24.5340023872, 32.9905601851, 68.5554944301, 69.1691724971, 37.3369520732, 52.3210070648, 66.9680225839, -0.823858069293};
test_label[2571] = '{69.1691724971};
test_output[2571] = '{0.502005999786};
############ END DEBUG ############*/
test_input[20576:20583] = '{32'h4010be62, 32'hc2ba6071, 32'hc2949f41, 32'h4227f348, 32'hc20ba96a, 32'hc19cf2d8, 32'hc250e406, 32'h4223f3d6};
test_label[2572] = '{32'hc2ba6071};
test_output[2572] = '{32'h43077d46};
/*############ DEBUG ############
test_input[20576:20583] = '{2.26162009405, -93.188359155, -74.3110427729, 41.9875795471, -34.9154434644, -19.6185768162, -52.2226775343, 40.9881215392};
test_label[2572] = '{-93.188359155};
test_output[2572] = '{135.489346183};
############ END DEBUG ############*/
test_input[20584:20591] = '{32'h413c5816, 32'h42b8a9d9, 32'h41e0d325, 32'hc29c4e8a, 32'hc2b5f5c3, 32'hc2b94600, 32'hc0cbe092, 32'h4211dc49};
test_label[2573] = '{32'h42b8a9d9};
test_output[2573] = '{32'h80000000};
/*############ DEBUG ############
test_input[20584:20591] = '{11.7715051271, 92.3317317489, 28.1030979067, -78.1533992844, -90.980001233, -92.6367220471, -6.37116333391, 36.4651224986};
test_label[2573] = '{92.3317317489};
test_output[2573] = '{-0.0};
############ END DEBUG ############*/
test_input[20592:20599] = '{32'h42c73bc3, 32'h41a82a61, 32'hc2615f3e, 32'hc27c29bf, 32'h42468fb9, 32'hc034da76, 32'h42b2b2f5, 32'h40069f4f};
test_label[2574] = '{32'hc2615f3e};
test_output[2574] = '{32'h431bf5b3};
/*############ DEBUG ############
test_input[20592:20599] = '{99.6167226218, 21.0206923128, -56.3430100668, -63.0407658991, 49.6403553774, -2.8258338043, 89.3495226682, 2.10347344886};
test_label[2574] = '{-56.3430100668};
test_output[2574] = '{155.959767443};
############ END DEBUG ############*/
test_input[20600:20607] = '{32'hc21ac1fb, 32'h41eefe83, 32'hc199c219, 32'hc2616674, 32'hc2503a4b, 32'hc2294050, 32'h428974f8, 32'hc204b022};
test_label[2575] = '{32'h428974f8};
test_output[2575] = '{32'h80000000};
/*############ DEBUG ############
test_input[20600:20607] = '{-38.6894352508, 29.874272919, -19.2197740233, -56.3500517103, -52.0569265859, -42.3128050345, 68.728457461, -33.1720064987};
test_label[2575] = '{68.728457461};
test_output[2575] = '{-0.0};
############ END DEBUG ############*/
test_input[20608:20615] = '{32'hc153ebd4, 32'h4287a466, 32'hc2c37e42, 32'hc294ca08, 32'hbfffb0b8, 32'hc08febea, 32'h421dc2f0, 32'h418233af};
test_label[2576] = '{32'hbfffb0b8};
test_output[2576] = '{32'h428ba329};
/*############ DEBUG ############
test_input[20608:20615] = '{-13.2450755628, 67.8210890104, -97.7465952509, -74.3945933611, -1.99758051073, -4.49754828329, 39.4403705595, 16.2752365248};
test_label[2576] = '{-1.99758051073};
test_output[2576] = '{69.8186695211};
############ END DEBUG ############*/
test_input[20616:20623] = '{32'hc16099a8, 32'h42c4ee12, 32'h40810aa8, 32'hc28ab260, 32'h41673778, 32'hc28fb053, 32'h424b376d, 32'h428d66eb};
test_label[2577] = '{32'h424b376d};
test_output[2577] = '{32'h423ea4b6};
/*############ DEBUG ############
test_input[20616:20623] = '{-14.0375139595, 98.46497862, 4.03255070827, -69.3483874438, 14.4510423188, -71.8443867372, 50.804127412, 70.7010080855};
test_label[2577] = '{50.804127412};
test_output[2577] = '{47.660851208};
############ END DEBUG ############*/
test_input[20624:20631] = '{32'h42a570c2, 32'hc0ff11ae, 32'h42b1f6d7, 32'h420f8a13, 32'hc26c6e48, 32'h424251ab, 32'hc2a68385, 32'h42c27ec9};
test_label[2578] = '{32'hc0ff11ae};
test_output[2578] = '{32'h42d27005};
/*############ DEBUG ############
test_input[20624:20631] = '{82.7202325833, -7.97090829594, 88.9821061096, 35.8848396461, -59.1076947812, 48.5797540668, -83.2568768558, 97.2476248398};
test_label[2578] = '{-7.97090829594};
test_output[2578] = '{105.218790829};
############ END DEBUG ############*/
test_input[20632:20639] = '{32'hc1df3abb, 32'hc250c480, 32'h42aa27ab, 32'hc24a9b3b, 32'hc2bfd022, 32'hc1106234, 32'hc2b95780, 32'hc29dbf30};
test_label[2579] = '{32'hc2b95780};
test_output[2579] = '{32'h4331bf95};
/*############ DEBUG ############
test_input[20632:20639] = '{-27.903676108, -52.1918957993, 85.0774727107, -50.6515936754, -95.9065069181, -9.02397495218, -92.6708956068, -78.8734138622};
test_label[2579] = '{-92.6708956068};
test_output[2579] = '{177.748368317};
############ END DEBUG ############*/
test_input[20640:20647] = '{32'hc1fd2efd, 32'h420afa35, 32'h424b3fbe, 32'hc1ae2d00, 32'h3d89ffd8, 32'h41759760, 32'h42488809, 32'hc252df59};
test_label[2580] = '{32'h424b3fbe};
test_output[2580] = '{32'h3ed1f473};
/*############ DEBUG ############
test_input[20640:20647] = '{-31.6479438445, 34.7443423297, 50.8122473746, -21.7719733062, 0.0673825130925, 15.3494567497, 50.1328459205, -52.718111343};
test_label[2580] = '{50.8122473746};
test_output[2580] = '{0.410068112551};
############ END DEBUG ############*/
test_input[20648:20655] = '{32'h413a5796, 32'hc2c56a79, 32'hc21854e7, 32'h42ac66a5, 32'h4280f05d, 32'hc27ed1d2, 32'h412bbe04, 32'hc180fa3e};
test_label[2581] = '{32'hc21854e7};
test_output[2581] = '{32'h42f89119};
/*############ DEBUG ############
test_input[20648:20655] = '{11.6463828377, -98.7079551127, -38.082911745, 86.2004792733, 64.4694617157, -63.7049021345, 10.7338909474, -16.1221894185};
test_label[2581] = '{-38.082911745};
test_output[2581] = '{124.283391019};
############ END DEBUG ############*/
test_input[20656:20663] = '{32'h4143f4b0, 32'hc1bc2041, 32'h4286d55c, 32'h424f471c, 32'h41fb9ce7, 32'hc02a5b07, 32'hc1f77a7c, 32'h419d4d51};
test_label[2582] = '{32'h41fb9ce7};
test_output[2582] = '{32'h420fdc45};
/*############ DEBUG ############
test_input[20656:20663] = '{12.2472383654, -23.5157491689, 67.4167184767, 51.8194414031, 31.4516115674, -2.66180596996, -30.9348069091, 19.662752152};
test_label[2582] = '{31.4516115674};
test_output[2582] = '{35.9651070776};
############ END DEBUG ############*/
test_input[20664:20671] = '{32'h42b4a66e, 32'hc0f168fb, 32'hc1eb8e64, 32'hc1aa514c, 32'h4256c98f, 32'hc1abf99d, 32'hc25760f9, 32'hc0344f9b};
test_label[2583] = '{32'h4256c98f};
test_output[2583] = '{32'h4212834e};
/*############ DEBUG ############
test_input[20664:20671] = '{90.3250608631, -7.54406503023, -29.4445260453, -21.2896949529, 53.6968350292, -21.4968808728, -53.8446985135, -2.81735882564};
test_label[2583] = '{53.6968350292};
test_output[2583] = '{36.6282258339};
############ END DEBUG ############*/
test_input[20672:20679] = '{32'h4144ef64, 32'hc22e290a, 32'hc22ce527, 32'hc1a62d24, 32'h4287a2a8, 32'hc2b4a278, 32'h429eefaf, 32'h40f92fca};
test_label[2584] = '{32'h4287a2a8};
test_output[2584] = '{32'h413a6844};
/*############ DEBUG ############
test_input[20672:20679] = '{12.3084448773, -43.5400762631, -43.2237828628, -20.7720420227, 67.8176869756, -90.3173226519, 79.4681341825, 7.78708361305};
test_label[2584] = '{67.8176869756};
test_output[2584] = '{11.650455922};
############ END DEBUG ############*/
test_input[20680:20687] = '{32'h40e0954a, 32'h4251a30b, 32'hc28b95ba, 32'hc1f9842f, 32'h429307ba, 32'h40b1e03c, 32'h4160b69d, 32'hc29fb1d7};
test_label[2585] = '{32'hc1f9842f};
test_output[2585] = '{32'h42d168c5};
/*############ DEBUG ############
test_input[20680:20687] = '{7.01822370132, 52.409222326, -69.7924342829, -31.1895420377, 73.5150894258, 5.55862258986, 14.0445834312, -79.8473419447};
test_label[2585] = '{-31.1895420377};
test_output[2585] = '{104.704631464};
############ END DEBUG ############*/
test_input[20688:20695] = '{32'h42a2cbd2, 32'hc2b656c7, 32'hc29625a7, 32'hc19810db, 32'hc2b5d631, 32'hc29c6f30, 32'h42137d19, 32'hc193adbf};
test_label[2586] = '{32'hc2b656c7};
test_output[2586] = '{32'h432c914c};
/*############ DEBUG ############
test_input[20688:20695] = '{81.3980831501, -91.1694893756, -75.0735367801, -19.0082302663, -90.9183456142, -78.21716547, 36.8721644079, -18.459836053};
test_label[2586] = '{-91.1694893756};
test_output[2586] = '{172.567572526};
############ END DEBUG ############*/
test_input[20696:20703] = '{32'h4115adc1, 32'h4236fb8a, 32'h429675df, 32'hc2bb5e46, 32'h42711e64, 32'hc213d154, 32'hc22877ae, 32'hc1bfe708};
test_label[2587] = '{32'hc22877ae};
test_output[2587] = '{32'h42eab1b6};
/*############ DEBUG ############
test_input[20696:20703] = '{9.35492027916, 45.7456441326, 75.2302156756, -93.6841276508, 60.2796782508, -36.9544207062, -42.11687505, -23.9878091577};
test_label[2587] = '{-42.11687505};
test_output[2587] = '{117.347091047};
############ END DEBUG ############*/
test_input[20704:20711] = '{32'h41dc7184, 32'hc1a9fb4a, 32'h41ff39bb, 32'h42c66675, 32'h425bbc66, 32'hc24ca3be, 32'hc21b93e0, 32'h4298c180};
test_label[2588] = '{32'hc21b93e0};
test_output[2588] = '{32'h430a1832};
/*############ DEBUG ############
test_input[20704:20711] = '{27.5554276565, -21.2476996346, 31.9031887884, 99.2001084549, 54.9339809721, -51.1599056014, -38.8944077641, 76.3779315939};
test_label[2588] = '{-38.8944077641};
test_output[2588] = '{138.094516219};
############ END DEBUG ############*/
test_input[20712:20719] = '{32'hc2a8dfe4, 32'h42baf92e, 32'hc2836481, 32'h41e18091, 32'h42a13f28, 32'h42b941c3, 32'h41c1a33f, 32'h427f2e9f};
test_label[2589] = '{32'h42a13f28};
test_output[2589] = '{32'h415377bd};
/*############ DEBUG ############
test_input[20712:20719] = '{-84.4372886543, 93.4866789469, -65.6962990448, 28.1877758513, 80.6233525509, 92.6284377008, 24.2047094906, 63.7955273739};
test_label[2589] = '{80.6233525509};
test_output[2589] = '{13.2167327003};
############ END DEBUG ############*/
test_input[20720:20727] = '{32'hc20ab727, 32'hc2633083, 32'hc161424f, 32'hc1def441, 32'h423cc22c, 32'h429ea672, 32'h41809bdd, 32'h4295fd27};
test_label[2590] = '{32'h423cc22c};
test_output[2590] = '{32'h4200981b};
/*############ DEBUG ############
test_input[20720:20727] = '{-34.6788614128, -56.7973733665, -14.0786882776, -27.869264561, 47.1896214261, 79.3250897101, 16.0761055091, 74.9944387923};
test_label[2590] = '{47.1896214261};
test_output[2590] = '{32.1485414361};
############ END DEBUG ############*/
test_input[20728:20735] = '{32'h41e9b32f, 32'hc23411cd, 32'hc247c0b3, 32'h427830ea, 32'h42813868, 32'h42b8ebc7, 32'h423f3b4f, 32'h42080bca};
test_label[2591] = '{32'h42813868};
test_output[2591] = '{32'h41decd7a};
/*############ DEBUG ############
test_input[20728:20735] = '{29.21249257, -45.0173824004, -49.9381822067, 62.0477671709, 64.6101690636, 92.4604997358, 47.8079167394, 34.0115120576};
test_label[2591] = '{64.6101690636};
test_output[2591] = '{27.8503306722};
############ END DEBUG ############*/
test_input[20736:20743] = '{32'hc01b2f9c, 32'h429a8b21, 32'h42847236, 32'hc18d83dd, 32'hc2c0dc04, 32'hc2b18536, 32'h429c7c9a, 32'h4111eeaa};
test_label[2592] = '{32'h4111eeaa};
test_output[2592] = '{32'h428ae31c};
/*############ DEBUG ############
test_input[20736:20743] = '{-2.4247807372, 77.2717327683, 66.2230697622, -17.689386685, -96.4297198928, -88.7601765743, 78.243360817, 9.12076723672};
test_label[2592] = '{9.12076723672};
test_output[2592] = '{69.4435695064};
############ END DEBUG ############*/
test_input[20744:20751] = '{32'hc2340d3e, 32'hc236f571, 32'hc227524d, 32'h416f8da3, 32'h423fcf58, 32'hc24e7524, 32'hc297dee9, 32'hc23de8b1};
test_label[2593] = '{32'h416f8da3};
test_output[2593] = '{32'h4203ebef};
/*############ DEBUG ############
test_input[20744:20751] = '{-45.0129329958, -45.739688687, -41.830373561, 14.9720794578, 47.9524850766, -51.6143962705, -75.9353701692, -47.4772361219};
test_label[2593] = '{14.9720794578};
test_output[2593] = '{32.9804056187};
############ END DEBUG ############*/
test_input[20752:20759] = '{32'hc1d3ef1b, 32'hc22c381e, 32'h42a31d35, 32'hc23bb9e1, 32'h42c70e44, 32'hc28eccf3, 32'hc2932a7f, 32'hc1ca5ce3};
test_label[2594] = '{32'hc22c381e};
test_output[2594] = '{32'h430e9529};
/*############ DEBUG ############
test_input[20752:20759] = '{-26.4917507311, -43.0548007206, 81.5570433919, -46.931521714, 99.5278620782, -71.4002937211, -73.583003147, -25.2953555142};
test_label[2594] = '{-43.0548007206};
test_output[2594] = '{142.582662814};
############ END DEBUG ############*/
test_input[20760:20767] = '{32'hc2a96d36, 32'h4116a7b8, 32'h422b7d70, 32'h415647e5, 32'hc057471d, 32'hc24be2bf, 32'h4282b749, 32'h42a9c299};
test_label[2595] = '{32'h422b7d70};
test_output[2595] = '{32'h422807c1};
/*############ DEBUG ############
test_input[20760:20767] = '{-84.713300314, 9.41594725577, 42.8724988686, 13.392552766, -3.36371548033, -50.971432748, 65.3579784325, 84.8800713552};
test_label[2595] = '{42.8724988686};
test_output[2595] = '{42.0075724899};
############ END DEBUG ############*/
test_input[20768:20775] = '{32'h3fc6b63e, 32'hc01efb90, 32'hc2b81c67, 32'h40fbdb0e, 32'h420faa9c, 32'h3dcdbdd4, 32'h4171ef87, 32'h41c03982};
test_label[2596] = '{32'h41c03982};
test_output[2596] = '{32'h413e3771};
/*############ DEBUG ############
test_input[20768:20775] = '{1.55243662009, -2.48410406189, -92.0554705745, 7.87049019124, 35.9166088773, 0.100459721926, 15.1209782677, 24.0280802329};
test_label[2596] = '{24.0280802329};
test_output[2596] = '{11.8885355141};
############ END DEBUG ############*/
test_input[20776:20783] = '{32'h41d4b86e, 32'hc2124df0, 32'h41d7f263, 32'hc2aed905, 32'hc28a2d65, 32'hc185665a, 32'hc2296a07, 32'hc2aca732};
test_label[2597] = '{32'hc185665a};
test_output[2597] = '{32'h4230b858};
/*############ DEBUG ############
test_input[20776:20783] = '{26.5900533903, -36.5761105197, 26.993353836, -87.4238686842, -69.0886604808, -16.6749762117, -42.3535425729, -86.3265534529};
test_label[2597] = '{-16.6749762117};
test_output[2597] = '{44.1800220988};
############ END DEBUG ############*/
test_input[20784:20791] = '{32'hc23d7a28, 32'hc28afaf0, 32'hc2b8d443, 32'h426e17f2, 32'hc268be58, 32'h428b47e8, 32'h42bf613f, 32'hc29d6b9f};
test_label[2598] = '{32'hc23d7a28};
test_output[2598] = '{32'h430f0f29};
/*############ DEBUG ############
test_input[20784:20791] = '{-47.3692914871, -69.4901117674, -92.4145720361, 59.523384864, -58.1858826565, 69.6404426961, 95.6899308647, -78.7102004256};
test_label[2598] = '{-47.3692914871};
test_output[2598] = '{143.059222352};
############ END DEBUG ############*/
test_input[20792:20799] = '{32'h420c34b1, 32'h424c0fe3, 32'hc1e0ddb0, 32'h4293c857, 32'hc200d053, 32'hc288abb9, 32'h420ded26, 32'h4253fa51};
test_label[2599] = '{32'hc288abb9};
test_output[2599] = '{32'h430e3a08};
/*############ DEBUG ############
test_input[20792:20799] = '{35.0514578461, 51.015513758, -28.1082466211, 73.8912873706, -32.2034410622, -68.335394123, 35.4815918687, 52.9944498153};
test_label[2599] = '{-68.335394123};
test_output[2599] = '{142.226681495};
############ END DEBUG ############*/
test_input[20800:20807] = '{32'h3f375822, 32'hc1fcf4bb, 32'h42af05e8, 32'hc28a4213, 32'h41ef82d5, 32'hc1872312, 32'hc24578f4, 32'hc295a01e};
test_label[2600] = '{32'hc1fcf4bb};
test_output[2600] = '{32'h42ee4316};
/*############ DEBUG ############
test_input[20800:20807] = '{0.716188570668, -31.6194966676, 87.511534258, -69.1290479218, 29.9388821027, -16.8921243028, -49.368120074, -74.812729488};
test_label[2600] = '{-31.6194966676};
test_output[2600] = '{119.131030926};
############ END DEBUG ############*/
test_input[20808:20815] = '{32'h41d6484a, 32'hc18d5785, 32'hc2878f1c, 32'h42c7cd1b, 32'hc20663d5, 32'hc249fd4e, 32'h411bb751, 32'hc1d9d488};
test_label[2601] = '{32'hc249fd4e};
test_output[2601] = '{32'h431665e1};
/*############ DEBUG ############
test_input[20808:20815] = '{26.7852979817, -17.6677349851, -67.7795134818, 99.9005933289, -33.597492464, -50.4973690827, 9.73225532033, -27.2287758398};
test_label[2601] = '{-50.4973690827};
test_output[2601] = '{150.397962412};
############ END DEBUG ############*/
test_input[20816:20823] = '{32'h41aa90b9, 32'hc257d776, 32'h42a27e45, 32'h4150280d, 32'hc18a7812, 32'hc2bb472f, 32'hc27e1f2a, 32'h41b0b55c};
test_label[2602] = '{32'hc18a7812};
test_output[2602] = '{32'h42c51c4a};
/*############ DEBUG ############
test_input[20816:20823] = '{21.3206651348, -53.9604126153, 81.2466231437, 13.0097784525, -17.3086272664, -93.6390332202, -63.5304344414, 22.0885543439};
test_label[2602] = '{-17.3086272664};
test_output[2602] = '{98.5552504101};
############ END DEBUG ############*/
test_input[20824:20831] = '{32'hc11f3f94, 32'hc14c5425, 32'h42007363, 32'hc29ef840, 32'hc2c15290, 32'hc1f72fd1, 32'h428ee125, 32'h42ad09af};
test_label[2603] = '{32'hc29ef840};
test_output[2603] = '{32'h432600f8};
/*############ DEBUG ############
test_input[20824:20831] = '{-9.9530217991, -12.7705426634, 32.1126827843, -79.4848668272, -96.6612543277, -30.8983470738, 71.4397337168, 86.5189099154};
test_label[2603] = '{-79.4848668272};
test_output[2603] = '{166.003777025};
############ END DEBUG ############*/
test_input[20832:20839] = '{32'h42c43928, 32'h4251e11e, 32'h42bc223c, 32'h42993810, 32'h4061e605, 32'hc2bc3bc7, 32'hc1f94935, 32'hc21bd32f};
test_label[2604] = '{32'hc1f94935};
test_output[2604] = '{32'h43014a2c};
/*############ DEBUG ############
test_input[20832:20839] = '{98.1116296521, 52.4698420441, 94.0668662744, 76.6094948215, 3.52966430644, -94.1167542027, -31.1607459556, -38.9562336887};
test_label[2604] = '{-31.1607459556};
test_output[2604] = '{129.289737856};
############ END DEBUG ############*/
test_input[20840:20847] = '{32'h42abfa8a, 32'h41de5997, 32'hc203004c, 32'h4255f027, 32'h425b51ea, 32'h410e6a2d, 32'h41b6bc89, 32'h429238a6};
test_label[2605] = '{32'h41de5997};
test_output[2605] = '{32'h4268c849};
/*############ DEBUG ############
test_input[20840:20847] = '{85.989333743, 27.7937452998, -32.7502898467, 53.4845247282, 54.829996096, 8.90092186187, 22.8420586521, 73.1106431213};
test_label[2605] = '{27.7937452998};
test_output[2605] = '{58.195590995};
############ END DEBUG ############*/
test_input[20848:20855] = '{32'hc0ee0bbe, 32'hc2154699, 32'h420859b5, 32'h42c0ffbc, 32'h4155b257, 32'hc21f2a31, 32'hc1bef611, 32'hc24d9355};
test_label[2606] = '{32'h420859b5};
test_output[2606] = '{32'h4279a5c3};
/*############ DEBUG ############
test_input[20848:20855] = '{-7.43893336226, -37.3189444408, 34.0876037507, 96.4994794238, 13.3560399234, -39.7912044255, -23.8701486717, -51.3938784799};
test_label[2606] = '{34.0876037507};
test_output[2606] = '{62.4118756731};
############ END DEBUG ############*/
test_input[20856:20863] = '{32'hc23839b4, 32'h428371ba, 32'h428cfc2c, 32'h41de3add, 32'h42998a02, 32'h429da84d, 32'hc25c46e4, 32'hc2468faa};
test_label[2607] = '{32'hc23839b4};
test_output[2607] = '{32'h42fa02bb};
/*############ DEBUG ############
test_input[20856:20863] = '{-46.0563488008, 65.7221189631, 70.4925247081, 27.7787416743, 76.7695458814, 78.8287113888, -55.0692291248, -49.6402985661};
test_label[2607] = '{-46.0563488008};
test_output[2607] = '{125.005330875};
############ END DEBUG ############*/
test_input[20864:20871] = '{32'hc28f427f, 32'hc1ee04a7, 32'hc282f22d, 32'h409a53ed, 32'h41927a02, 32'h41b1ae66, 32'hc2b8ee2b, 32'h4233dfe3};
test_label[2608] = '{32'h4233dfe3};
test_output[2608] = '{32'h2f128f30};
/*############ DEBUG ############
test_input[20864:20871] = '{-71.6298737679, -29.7522720481, -65.4729994086, 4.82274496664, 18.3095736343, 22.2101547525, -92.4651711817, 44.9686397925};
test_label[2608] = '{44.9686397925};
test_output[2608] = '{1.33294930658e-10};
############ END DEBUG ############*/
test_input[20872:20879] = '{32'hc1453037, 32'hc2099881, 32'hc2937e1e, 32'hc26e18f2, 32'hc298db34, 32'hc28e3d0f, 32'hc25866f3, 32'hc0c5f0a7};
test_label[2609] = '{32'hc298db34};
test_output[2609] = '{32'h428c7d44};
/*############ DEBUG ############
test_input[20872:20879] = '{-12.3242708484, -34.3989283389, -73.7463201822, -59.5243595107, -76.4281285482, -71.119257802, -54.1005373289, -6.18562641471};
test_label[2609] = '{-76.4281285482};
test_output[2609] = '{70.2446576554};
############ END DEBUG ############*/
test_input[20880:20887] = '{32'hc1d7655f, 32'hc28fdb48, 32'hc2b1a802, 32'h42935b02, 32'hc2999c75, 32'hc08d9706, 32'hc2305038, 32'h42161a1d};
test_label[2610] = '{32'hc28fdb48};
test_output[2610] = '{32'h43119b25};
/*############ DEBUG ############
test_input[20880:20887] = '{-26.9244982683, -71.9282815038, -88.8281374895, 73.677751259, -76.8055784158, -4.42468559268, -44.0783395438, 37.5255018646};
test_label[2610] = '{-71.9282815038};
test_output[2610] = '{145.606032763};
############ END DEBUG ############*/
test_input[20888:20895] = '{32'h41a87d0d, 32'h42257a42, 32'h427e4c9e, 32'h41932cc0, 32'h41536dc9, 32'hc27b4083, 32'hc21f822b, 32'hc2a005b5};
test_label[2611] = '{32'h41536dc9};
test_output[2611] = '{32'h4249712b};
/*############ DEBUG ############
test_input[20888:20895] = '{21.0610597328, 41.369391144, 63.5748197388, 18.396850108, 13.2143028303, -62.8129998656, -39.8771158812, -80.0111443671};
test_label[2611] = '{13.2143028303};
test_output[2611] = '{50.3605169087};
############ END DEBUG ############*/
test_input[20896:20903] = '{32'h41f478ac, 32'hc28ae564, 32'h4148b43f, 32'h41a75dc5, 32'h3fe327d5, 32'h42825191, 32'h42a5c1f0, 32'hc107ad64};
test_label[2612] = '{32'h4148b43f};
test_output[2612] = '{32'h428cab68};
/*############ DEBUG ############
test_input[20896:20903] = '{30.558922358, -69.448029445, 12.5440049964, 20.9207851941, 1.77465312914, 65.1593062118, 82.8787827881, -8.47983177912};
test_label[2612] = '{12.5440049964};
test_output[2612] = '{70.3347778119};
############ END DEBUG ############*/
test_input[20904:20911] = '{32'h421f3ea5, 32'hc2bdf8cd, 32'h42095b94, 32'h42405de5, 32'h429823c6, 32'h417ca355, 32'h418ee21b, 32'hc12f4989};
test_label[2613] = '{32'hc2bdf8cd};
test_output[2613] = '{32'h432b0e4a};
/*############ DEBUG ############
test_input[20904:20911] = '{39.8111773992, -94.9859383216, 34.3394329896, 48.0916921167, 76.0698735917, 15.7898756991, 17.8604035018, -10.9554524792};
test_label[2613] = '{-94.9859383216};
test_output[2613] = '{171.055811913};
############ END DEBUG ############*/
test_input[20912:20919] = '{32'hc02d68b7, 32'h421c019d, 32'h427c4dfc, 32'h424cc376, 32'hc2a29a68, 32'hc1fdb848, 32'h427b6039, 32'h4297183d};
test_label[2614] = '{32'hc2a29a68};
test_output[2614] = '{32'h431cd953};
/*############ DEBUG ############
test_input[20912:20919] = '{-2.70951634346, 39.0015771332, 63.0761579143, 51.1908793589, -81.3015773859, -31.7149817039, 62.8439680075, 75.5473433008};
test_label[2614] = '{-81.3015773859};
test_output[2614] = '{156.848927563};
############ END DEBUG ############*/
test_input[20920:20927] = '{32'hc25679bd, 32'h421a5685, 32'h429412ca, 32'hc1fae8a5, 32'hc24afcfe, 32'hc2c52489, 32'h428f0f8e, 32'hc298ec11};
test_label[2615] = '{32'h421a5685};
test_output[2615] = '{32'h420e1f5a};
/*############ DEBUG ############
test_input[20920:20927] = '{-53.6188844172, 38.584491224, 74.0366979219, -31.3635954349, -50.747064213, -98.5713605422, 71.5303813238, -76.4610654479};
test_label[2615] = '{38.584491224};
test_output[2615] = '{35.5306186625};
############ END DEBUG ############*/
test_input[20928:20935] = '{32'hc2c5b88c, 32'hc24cf429, 32'h42a30c7a, 32'h42ae37a8, 32'hc1df7dcc, 32'h425da2aa, 32'hc2c52f91, 32'h416aa453};
test_label[2616] = '{32'h425da2aa};
test_output[2616] = '{32'h41fda0f8};
/*############ DEBUG ############
test_input[20928:20935] = '{-98.8604400775, -51.2384359565, 81.5243698993, 87.1087018887, -27.9364251536, 55.4088523563, -98.592906337, 14.6651183848};
test_label[2616] = '{55.4088523563};
test_output[2616] = '{31.7035987535};
############ END DEBUG ############*/
test_input[20936:20943] = '{32'hc28d92c6, 32'hc253062a, 32'hc2569bd8, 32'hc2049fe5, 32'h41ca9412, 32'h41f338a9, 32'hc258cf42, 32'h426fb584};
test_label[2617] = '{32'hc2049fe5};
test_output[2617] = '{32'h42ba2ab5};
/*############ DEBUG ############
test_input[20936:20943] = '{-70.7866700192, -52.756021199, -53.6521926866, -33.1561477147, 25.3222992813, 30.4026666149, -54.2024019454, 59.9272628265};
test_label[2617] = '{-33.1561477147};
test_output[2617] = '{93.0834105413};
############ END DEBUG ############*/
test_input[20944:20951] = '{32'h4229da92, 32'hc22a61b3, 32'h421ab836, 32'hc1bb679a, 32'hc273f149, 32'h416ea829, 32'hc2a7cab3, 32'hc201b55b};
test_label[2618] = '{32'hc273f149};
test_output[2618] = '{32'h42cef171};
/*############ DEBUG ############
test_input[20944:20951] = '{42.4634459849, -42.5954112413, 38.6798924873, -23.4255872807, -60.9856311423, 14.9160543382, -83.8958960685, -32.4271063879};
test_label[2618] = '{-60.9856311423};
test_output[2618] = '{103.471564124};
############ END DEBUG ############*/
test_input[20952:20959] = '{32'hc2ae3eaf, 32'hc282e9e9, 32'h42b6fa0b, 32'h416be26d, 32'hc08be167, 32'h42a73a88, 32'h4291dfbc, 32'h422620a7};
test_label[2619] = '{32'h42b6fa0b};
test_output[2619] = '{32'h39c773ec};
/*############ DEBUG ############
test_input[20952:20959] = '{-87.1224283305, -65.4568526686, 91.4883684365, 14.7427799182, -4.37126505065, 83.6143168432, 72.9369827756, 41.5318880541};
test_label[2619] = '{91.4883684365};
test_output[2619] = '{0.000380426049332};
############ END DEBUG ############*/
test_input[20960:20967] = '{32'h42a1aef2, 32'h41fd80ab, 32'hc2bf133e, 32'hc291d64a, 32'hc191f202, 32'hc220d472, 32'hbf8139a6, 32'hc2a4c37c};
test_label[2620] = '{32'hc191f202};
test_output[2620] = '{32'h42c62b72};
/*############ DEBUG ############
test_input[20960:20967] = '{80.8416886194, 31.6878262179, -95.5375859019, -72.9185342367, -18.2431671887, -40.2074661449, -1.0095718308, -82.3818085075};
test_label[2620] = '{-18.2431671887};
test_output[2620] = '{99.0848558082};
############ END DEBUG ############*/
test_input[20968:20975] = '{32'h412371b4, 32'h40ced822, 32'hc1775519, 32'h42411189, 32'hc25b35a2, 32'hc1712450, 32'h42c26e6f, 32'h42754a0f};
test_label[2621] = '{32'h412371b4};
test_output[2621] = '{32'h42ae0039};
/*############ DEBUG ############
test_input[20968:20975] = '{10.215259902, 6.46388338402, -15.4582762016, 48.2671239279, -54.8023747909, -15.071365772, 97.2156912579, 61.3223238392};
test_label[2621] = '{10.215259902};
test_output[2621] = '{87.0004313559};
############ END DEBUG ############*/
test_input[20976:20983] = '{32'hc2601dab, 32'h42a08648, 32'h429add3b, 32'h4246c4e2, 32'h41fff29f, 32'hc25110d8, 32'hc1ebe4b2, 32'h428110f7};
test_label[2622] = '{32'hc25110d8};
test_output[2622] = '{32'h43049607};
/*############ DEBUG ############
test_input[20976:20983] = '{-56.0289742321, 80.2622649794, 77.4320906763, 49.692270027, 31.9934664712, -52.2664484421, -29.4866674979, 64.5331312805};
test_label[2622] = '{-52.2664484421};
test_output[2622] = '{132.586041053};
############ END DEBUG ############*/
test_input[20984:20991] = '{32'hc282c491, 32'hc114c9f4, 32'hc2992af6, 32'h4253a63f, 32'hc2ad32fb, 32'h4203320d, 32'h4282d3b4, 32'h42217079};
test_label[2623] = '{32'h4282d3b4};
test_output[2623] = '{32'h3679cf2b};
/*############ DEBUG ############
test_input[20984:20991] = '{-65.3839162131, -9.29930450944, -76.5839079562, 52.9123500519, -86.5995732631, 32.798878005, 65.4134807799, 40.3598347265};
test_label[2623] = '{65.4134807799};
test_output[2623] = '{3.7224479636e-06};
############ END DEBUG ############*/
test_input[20992:20999] = '{32'h423278ac, 32'h4174198b, 32'h4289745e, 32'h416bcd50, 32'h4245d095, 32'h428fdd11, 32'h429456ba, 32'h419660ed};
test_label[2624] = '{32'h416bcd50};
test_output[2624] = '{32'h426e25f3};
/*############ DEBUG ############
test_input[20992:20999] = '{44.6178448034, 15.2562361724, 68.727279632, 14.7376247263, 49.4536947532, 71.9317667826, 74.1693870773, 18.7973277638};
test_label[2624] = '{14.7376247263};
test_output[2624] = '{59.537061109};
############ END DEBUG ############*/
test_input[21000:21007] = '{32'hc20da8b7, 32'hc1cb890d, 32'hc253a25e, 32'hc2972b17, 32'hc181474d, 32'h4092311e, 32'hc1b95e0f, 32'hc2a42270};
test_label[2625] = '{32'hc2972b17};
test_output[2625] = '{32'h42a04e29};
/*############ DEBUG ############
test_input[21000:21007] = '{-35.414758898, -25.4419184599, -52.9085625475, -75.5841592181, -16.1598142087, 4.56849574604, -23.1709274196, -82.0672635007};
test_label[2625] = '{-75.5841592181};
test_output[2625] = '{80.1526549652};
############ END DEBUG ############*/
test_input[21008:21015] = '{32'h4217ddd9, 32'hc2b9d28e, 32'h4138a65b, 32'hc2bb450f, 32'hc23a03c1, 32'hc2b1e23f, 32'h424ae8ac, 32'hc2aec638};
test_label[2626] = '{32'h4138a65b};
test_output[2626] = '{32'h421cbf17};
/*############ DEBUG ############
test_input[21008:21015] = '{37.9666462978, -92.9112432504, 11.5406138941, -93.6348796671, -46.5036660225, -88.9418862597, 50.7272204052, -87.3871460243};
test_label[2626] = '{11.5406138941};
test_output[2626] = '{39.1866093828};
############ END DEBUG ############*/
test_input[21016:21023] = '{32'hc2850499, 32'h41159a55, 32'hc2b7bfa1, 32'h4294607e, 32'hc29ddc36, 32'hc26b8371, 32'hc2350bbe, 32'h410ae0ec};
test_label[2627] = '{32'h410ae0ec};
test_output[2627] = '{32'h42830460};
/*############ DEBUG ############
test_input[21016:21023] = '{-66.5089770442, 9.35017906809, -91.8742755307, 74.1884584772, -78.9301008777, -58.8783597632, -45.2614655976, 8.67991259669};
test_label[2627] = '{8.67991259669};
test_output[2627] = '{65.5085458805};
############ END DEBUG ############*/
test_input[21024:21031] = '{32'hc2a21659, 32'hc2acb540, 32'hc2bb372f, 32'h42994933, 32'hc29f2372, 32'hc1882a51, 32'hc26e2639, 32'h429c177c};
test_label[2628] = '{32'hc26e2639};
test_output[2628] = '{32'h4309cd94};
/*############ DEBUG ############
test_input[21024:21031] = '{-81.0436469729, -86.3540020385, -93.6077779233, 76.6429637349, -79.5692302559, -17.0206627755, -59.5373285815, 78.0458648313};
test_label[2628] = '{-59.5373285815};
test_output[2628] = '{137.803037606};
############ END DEBUG ############*/
test_input[21032:21039] = '{32'hc0da8cee, 32'hc2b42a62, 32'hc29f0faf, 32'hc2a487e9, 32'h42b72c2f, 32'h428a262e, 32'hc1c9baca, 32'hc1747689};
test_label[2629] = '{32'hc0da8cee};
test_output[2629] = '{32'h42c4d4fe};
/*############ DEBUG ############
test_input[21032:21039] = '{-6.82970315942, -90.0827815884, -79.5306292243, -82.2654491505, 91.5862944198, 69.0745726023, -25.2162047294, -15.2789390804};
test_label[2629] = '{-6.82970315942};
test_output[2629] = '{98.4159975794};
############ END DEBUG ############*/
test_input[21040:21047] = '{32'h428efb0f, 32'hc2c1b071, 32'hc2ba3fa8, 32'h42c27542, 32'h420f374b, 32'h42c369f2, 32'h42ad743c, 32'h41e17089};
test_label[2630] = '{32'h42c369f2};
test_output[2630] = '{32'h3ef708b3};
/*############ DEBUG ############
test_input[21040:21047] = '{71.4903511167, -96.8446118903, -93.1243250569, 97.2290196964, 35.8039984038, 97.706920731, 86.727019056, 28.1799482487};
test_label[2630] = '{97.706920731};
test_output[2630] = '{0.482488247055};
############ END DEBUG ############*/
test_input[21048:21055] = '{32'h42808c9b, 32'h42c58e22, 32'h4296142d, 32'h429f414c, 32'hc27f97c9, 32'hc262d545, 32'h4228246a, 32'h42898e4f};
test_label[2631] = '{32'hc27f97c9};
test_output[2631] = '{32'h4322ad03};
/*############ DEBUG ############
test_input[21048:21055] = '{64.2746195438, 98.777603658, 75.0394088994, 79.6275315041, -63.8982267692, -56.7082699579, 42.0355596693, 68.7779438878};
test_label[2631] = '{-63.8982267692};
test_output[2631] = '{162.675830432};
############ END DEBUG ############*/
test_input[21056:21063] = '{32'hc163f4a2, 32'h428fac89, 32'h42c370a3, 32'hc0ba56a2, 32'h400cb4c7, 32'hc2ae12bc, 32'hc287bb2f, 32'hc2324723};
test_label[2632] = '{32'h428fac89};
test_output[2632] = '{32'h41cf1066};
/*############ DEBUG ############
test_input[21056:21063] = '{-14.2472252408, 71.8369857501, 97.7199933324, -5.82307509951, 2.19853386965, -87.0365886405, -67.8655915899, -44.5694677593};
test_label[2632] = '{71.8369857501};
test_output[2632] = '{25.8830075823};
############ END DEBUG ############*/
test_input[21064:21071] = '{32'h41d49e15, 32'hc2bb1858, 32'h42b772c9, 32'h42b34889, 32'hc28b80f4, 32'hc2aae1af, 32'hc28cf544, 32'h41b02d85};
test_label[2633] = '{32'h42b772c9};
test_output[2633] = '{32'h3df08529};
/*############ DEBUG ############
test_input[21064:21071] = '{26.5771889239, -93.5475436259, 91.7241892826, 89.6416695658, -69.7518590365, -85.4407884808, -70.479036483, 22.0222265836};
test_label[2633] = '{91.7241892826};
test_output[2633] = '{0.117441483734};
############ END DEBUG ############*/
test_input[21072:21079] = '{32'hc1e1afbc, 32'h4299495c, 32'hc1a91bc3, 32'h41d48010, 32'h426752bf, 32'h42c7029b, 32'hc055e344, 32'h42a29008};
test_label[2634] = '{32'h42a29008};
test_output[2634] = '{32'h4191ca4c};
/*############ DEBUG ############
test_input[21072:21079] = '{-28.2108086092, 76.6432778645, -21.1385547345, 26.5625311616, 57.830808173, 99.5050871545, -3.34199608679, 81.2813086052};
test_label[2634] = '{81.2813086052};
test_output[2634] = '{18.2237785615};
############ END DEBUG ############*/
test_input[21080:21087] = '{32'hc2c7acc2, 32'h42bf8946, 32'hc297b829, 32'hc1e02474, 32'h42157003, 32'hc2951fb6, 32'h4187801b, 32'h42ba0045};
test_label[2635] = '{32'h42ba0045};
test_output[2635] = '{32'h40350625};
/*############ DEBUG ############
test_input[21080:21087] = '{-99.8374141182, 95.7681093426, -75.8596875317, -28.0177984257, 37.359386845, -74.5619358032, 16.9375507128, 93.0005291266};
test_label[2635] = '{93.0005291266};
test_output[2635] = '{2.82850015122};
############ END DEBUG ############*/
test_input[21088:21095] = '{32'h419663c2, 32'hc2108a70, 32'hc24eeadc, 32'hc250f3de, 32'hc0d48830, 32'h42a97e26, 32'h4222c03d, 32'h419dc868};
test_label[2636] = '{32'h42a97e26};
test_output[2636] = '{32'h80000000};
/*############ DEBUG ############
test_input[21088:21095] = '{18.7987096008, -36.1351929097, -51.7293531765, -52.2381518493, -6.64162448449, 84.7463853278, 40.6877330831, 19.7228542688};
test_label[2636] = '{84.7463853278};
test_output[2636] = '{-0.0};
############ END DEBUG ############*/
test_input[21096:21103] = '{32'hc2200ce9, 32'h429716cf, 32'h4039d3dc, 32'h42aff01d, 32'hc0bb50f6, 32'hc2b72f0e, 32'h429c1278, 32'h42314926};
test_label[2637] = '{32'h42aff01d};
test_output[2637] = '{32'h385c7ce9};
/*############ DEBUG ############
test_input[21096:21103] = '{-40.0126079287, 75.5445448125, 2.90355577186, 87.9689736437, -5.85363292296, -91.5919068537, 78.0360697868, 44.3214322181};
test_label[2637] = '{87.9689736437};
test_output[2637] = '{5.25684208182e-05};
############ END DEBUG ############*/
test_input[21104:21111] = '{32'h4156edc7, 32'h4200ac22, 32'hc1d2dca0, 32'hc2491a5f, 32'h42505579, 32'hc028ce78, 32'hc29088f4, 32'hc19e998b};
test_label[2638] = '{32'h4200ac22};
test_output[2638] = '{32'h419f52af};
/*############ DEBUG ############
test_input[21104:21111] = '{13.4330511056, 32.1680991237, -26.3577279354, -50.2757534005, 52.0834712631, -2.63760196287, -72.2674876693, -19.8249714517};
test_label[2638] = '{32.1680991237};
test_output[2638] = '{19.9153721417};
############ END DEBUG ############*/
test_input[21112:21119] = '{32'h4263a1b8, 32'hc22438cf, 32'h42c424e5, 32'h41bc458d, 32'h42959d25, 32'hc1ab1314, 32'hc294765e, 32'h421ee163};
test_label[2639] = '{32'hc22438cf};
test_output[2639] = '{32'h430b20a6};
/*############ DEBUG ############
test_input[21112:21119] = '{56.9079275385, -41.055477852, 98.0720593023, 23.5339598464, 74.8069246604, -21.3843153152, -74.2311832237, 39.720102401};
test_label[2639] = '{-41.055477852};
test_output[2639] = '{139.127537154};
############ END DEBUG ############*/
test_input[21120:21127] = '{32'h4164a587, 32'hc1e4b6b2, 32'h42ab7243, 32'h42197969, 32'h42344983, 32'h4195abac, 32'hc0effba7, 32'hc2c59d67};
test_label[2640] = '{32'h42197969};
test_output[2640] = '{32'h423d6b1d};
/*############ DEBUG ############
test_input[21120:21127] = '{14.2904120398, -28.5892073306, 85.7231667042, 38.3685643139, 45.0717877414, 18.7088242782, -7.4994690461, -98.8074251739};
test_label[2640] = '{38.3685643139};
test_output[2640] = '{47.3546023904};
############ END DEBUG ############*/
test_input[21128:21135] = '{32'h42ace995, 32'h40a2b639, 32'hc1aa5cb3, 32'h41b5fd1e, 32'hc1b8a8d3, 32'hc06271ce, 32'hc29460ee, 32'h41f67c11};
test_label[2641] = '{32'h40a2b639};
test_output[2641] = '{32'h42a2be32};
/*############ DEBUG ############
test_input[21128:21135] = '{86.4562159675, 5.08474396944, -21.2952624941, 22.7485923562, -23.0824336385, -3.53819610506, -74.1893137147, 30.8105788022};
test_label[2641] = '{5.08474396944};
test_output[2641] = '{81.3714719981};
############ END DEBUG ############*/
test_input[21136:21143] = '{32'hc23d621e, 32'hc295d522, 32'h42a9625c, 32'hc1c1a7f7, 32'hc2b0f211, 32'h421c73b6, 32'h424b5794, 32'hc2634438};
test_label[2642] = '{32'hc2b0f211};
test_output[2642] = '{32'h432d2a36};
/*############ DEBUG ############
test_input[21136:21143] = '{-47.345818572, -74.9162727912, 84.6921056424, -24.2070140178, -88.4727835474, 39.112999541, 50.835527288, -56.8166192587};
test_label[2642] = '{-88.4727835474};
test_output[2642] = '{173.16488919};
############ END DEBUG ############*/
test_input[21144:21151] = '{32'h42abd3a4, 32'hc23f1a28, 32'h421e4da3, 32'hc1ab8f25, 32'h419676b2, 32'h421eca23, 32'h42b03b5d, 32'hc243f9cf};
test_label[2643] = '{32'h421eca23};
test_output[2643] = '{32'h424217ed};
/*############ DEBUG ############
test_input[21144:21151] = '{85.9133614918, -47.7755442456, 39.5758167218, -21.4448955646, 18.8079572405, 39.6974006006, 88.1159407519, -48.9939547865};
test_label[2643] = '{39.6974006006};
test_output[2643] = '{48.5233664871};
############ END DEBUG ############*/
test_input[21152:21159] = '{32'h42c70c97, 32'h4291e985, 32'hc290f9bb, 32'h41f831dc, 32'hc1d15943, 32'hc12dd376, 32'h41f1c936, 32'hc287b4fe};
test_label[2644] = '{32'hc12dd376};
test_output[2644] = '{32'h42dcc705};
/*############ DEBUG ############
test_input[21152:21159] = '{99.5245875749, 72.9560916528, -72.4877546447, 31.0243455159, -26.168585409, -10.8641259706, 30.2232476222, -67.8535026562};
test_label[2644] = '{-10.8641259706};
test_output[2644] = '{110.388713545};
############ END DEBUG ############*/
test_input[21160:21167] = '{32'hc10b3369, 32'hc0bb19da, 32'hc203840e, 32'h426dc06d, 32'h41433706, 32'h429ae83c, 32'h421687de, 32'h420b73c2};
test_label[2645] = '{32'h429ae83c};
test_output[2645] = '{32'h3280caa2};
/*############ DEBUG ############
test_input[21160:21167] = '{-8.70005092144, -5.84690571725, -32.8789583946, 59.437917567, 12.200933076, 77.4535794741, 37.6326843477, 34.8630429926};
test_label[2645] = '{77.4535794741};
test_output[2645] = '{1.49933073748e-08};
############ END DEBUG ############*/
test_input[21168:21175] = '{32'h42ad3ff6, 32'h427abd2d, 32'h429ed134, 32'hc2acaa56, 32'h426ce3f4, 32'hc2c4f4fe, 32'h4232b18c, 32'hc29d7842};
test_label[2646] = '{32'h4232b18c};
test_output[2646] = '{32'h4227cf1f};
/*############ DEBUG ############
test_input[21168:21175] = '{86.6249208584, 62.6847421012, 79.4085993985, -86.3326863509, 59.2226107784, -98.4785002159, 44.6733872487, -78.7348777142};
test_label[2646] = '{44.6733872487};
test_output[2646] = '{41.9522678395};
############ END DEBUG ############*/
test_input[21176:21183] = '{32'h412b930e, 32'h427ba967, 32'hc19e71ee, 32'hc25e1d85, 32'hc100167b, 32'hc218f70c, 32'hc26251bd, 32'hc1a4e18e};
test_label[2647] = '{32'hc26251bd};
test_output[2647] = '{32'h42eefd92};
/*############ DEBUG ############
test_input[21176:21183] = '{10.7234017209, 62.915431035, -19.8056297082, -55.5288272205, -8.00548861262, -38.2412561444, -56.5798233009, -20.6101338057};
test_label[2647] = '{-56.5798233009};
test_output[2647] = '{119.495254336};
############ END DEBUG ############*/
test_input[21184:21191] = '{32'hc24eb1fc, 32'hc264dffd, 32'hc1c4f6b0, 32'h42b6f3aa, 32'hc121efe2, 32'h4237ec27, 32'h4167a42e, 32'h42321943};
test_label[2648] = '{32'h4237ec27};
test_output[2648] = '{32'h4235fb2d};
/*############ DEBUG ############
test_input[21184:21191] = '{-51.6738114565, -57.2187370434, -24.6204525186, 91.4759061758, -10.1210649616, 45.9806175285, 14.4775824729, 44.5246694021};
test_label[2648] = '{45.9806175285};
test_output[2648] = '{45.4952886473};
############ END DEBUG ############*/
test_input[21192:21199] = '{32'hc1b938b3, 32'h425e56df, 32'hc111dd50, 32'hc2befdde, 32'h42857d12, 32'hc2a5329b, 32'h424c3acf, 32'h42aba98f};
test_label[2649] = '{32'hc2befdde};
test_output[2649] = '{32'h433553b6};
/*############ DEBUG ############
test_input[21192:21199] = '{-23.1526846104, 55.584835291, -9.11653102276, -95.4958322572, 66.7442803467, -82.5988366581, 51.0574298257, 85.8311661303};
test_label[2649] = '{-95.4958322572};
test_output[2649] = '{181.326998393};
############ END DEBUG ############*/
test_input[21200:21207] = '{32'h42c3a67f, 32'hc29f070a, 32'hc277a704, 32'hc2863b63, 32'h423ee0a7, 32'h42851776, 32'h416a4444, 32'h4258335d};
test_label[2650] = '{32'h42851776};
test_output[2650] = '{32'h41fa3c27};
/*############ DEBUG ############
test_input[21200:21207] = '{97.825191015, -79.5137496437, -61.9131016123, -67.1159917232, 47.7193851676, 66.5458194409, 14.6416667565, 54.050159172};
test_label[2650] = '{66.5458194409};
test_output[2650] = '{31.2793715742};
############ END DEBUG ############*/
test_input[21208:21215] = '{32'h429e2a60, 32'hc0b7b89f, 32'hc21846b0, 32'hc20a5a7e, 32'h427369da, 32'h42b310c6, 32'h42498726, 32'hc2524aaf};
test_label[2651] = '{32'h427369da};
test_output[2651] = '{32'h41e56f73};
/*############ DEBUG ############
test_input[21208:21215] = '{79.0827666779, -5.74128679876, -38.069029056, -34.588371484, 60.8533703595, 89.5327596482, 50.3819820782, -52.5729321326};
test_label[2651] = '{60.8533703595};
test_output[2651] = '{28.6794182367};
############ END DEBUG ############*/
test_input[21216:21223] = '{32'hc097db5f, 32'h42a1cb72, 32'h42155aee, 32'hc28aae52, 32'h41c668b1, 32'hc25ab7d3, 32'hc24259c6, 32'hc2944aad};
test_label[2652] = '{32'hc24259c6};
test_output[2652] = '{32'h43017c2b};
/*############ DEBUG ############
test_input[21216:21223] = '{-4.745528708, 80.8973540596, 37.3387977294, -69.3404722043, 24.8011194384, -54.6795159135, -48.5876699941, -74.1458477232};
test_label[2652] = '{-48.5876699941};
test_output[2652] = '{129.485024054};
############ END DEBUG ############*/
test_input[21224:21231] = '{32'h41ad5468, 32'hc21c7ff0, 32'h42bab386, 32'h3f5ff60c, 32'h427cc82b, 32'hc0bac944, 32'hc2a9a107, 32'hc202fdeb};
test_label[2653] = '{32'hc202fdeb};
test_output[2653] = '{32'h42fc327c};
/*############ DEBUG ############
test_input[21224:21231] = '{21.6662135534, -39.1249387256, 93.3506328388, 0.874848140537, 63.1954783647, -5.83706832374, -84.8145053825, -32.7479670134};
test_label[2653] = '{-32.7479670134};
test_output[2653] = '{126.098599852};
############ END DEBUG ############*/
test_input[21232:21239] = '{32'hbe8048f7, 32'hbe823917, 32'h428141ba, 32'h41f56d0e, 32'hc2b7bfa9, 32'h41907120, 32'hc2bd2c80, 32'hc0c9ef0c};
test_label[2654] = '{32'hc2bd2c80};
test_output[2654] = '{32'h431f371d};
/*############ DEBUG ############
test_input[21232:21239] = '{-0.250556683782, -0.2543418037, 64.6283741864, 30.6782489669, -91.8743370005, 18.0552368362, -94.5869114363, -6.31043053319};
test_label[2654] = '{-94.5869114363};
test_output[2654] = '{159.215285623};
############ END DEBUG ############*/
test_input[21240:21247] = '{32'h4297098c, 32'hc1b2daa8, 32'h417a1363, 32'h42b28b1c, 32'h4295b8d4, 32'h4282afed, 32'h425fcb52, 32'hc1228fac};
test_label[2655] = '{32'h4295b8d4};
test_output[2655] = '{32'h41669248};
/*############ DEBUG ############
test_input[21240:21247] = '{75.5186459425, -22.3567660043, 15.6297326842, 89.2717002644, 74.8609891359, 65.3436069223, 55.9485540272, -10.1600764899};
test_label[2655] = '{74.8609891359};
test_output[2655] = '{14.4107127445};
############ END DEBUG ############*/
test_input[21248:21255] = '{32'h42b4ab1b, 32'hc27ff3c2, 32'h42bc0585, 32'hc19c387a, 32'hc19efea7, 32'h42048d21, 32'hc18ebba4, 32'h415ed6cf};
test_label[2656] = '{32'h415ed6cf};
test_output[2656] = '{32'h42a03778};
/*############ DEBUG ############
test_input[21248:21255] = '{90.3341929925, -63.9880456636, 94.010783325, -19.5275770673, -19.8743428028, 33.1378192936, -17.8416215148, 13.9274431792};
test_label[2656] = '{13.9274431792};
test_output[2656] = '{80.108334297};
############ END DEBUG ############*/
test_input[21256:21263] = '{32'h42822d23, 32'h419ea7b5, 32'hc24794d3, 32'h41dc1d71, 32'hc21e91cf, 32'hc28b914f, 32'hc2973904, 32'h4248affc};
test_label[2657] = '{32'h4248affc};
test_output[2657] = '{32'h416ea929};
/*############ DEBUG ############
test_input[21256:21263] = '{65.088156808, 19.83188832, -49.8953356326, 27.51437664, -39.6423921382, -69.7838054705, -75.6113555849, 50.1718584445};
test_label[2657] = '{50.1718584445};
test_output[2657] = '{14.9162986962};
############ END DEBUG ############*/
test_input[21264:21271] = '{32'h41f79dd3, 32'h423bfa1d, 32'h42937dba, 32'hc283a0c2, 32'hc29a3162, 32'h413067a5, 32'h42c089f7, 32'hc26d2593};
test_label[2658] = '{32'h413067a5};
test_output[2658] = '{32'h42aa7d02};
/*############ DEBUG ############
test_input[21264:21271] = '{30.9520632654, 46.9942517582, 73.7455612739, -65.8139809116, -77.0964473873, 11.0253036821, 96.2694618643, -59.2866934879};
test_label[2658] = '{11.0253036821};
test_output[2658] = '{85.2441581824};
############ END DEBUG ############*/
test_input[21272:21279] = '{32'h428b0da6, 32'hc2b4ae8e, 32'hc2ada806, 32'hc1279670, 32'hc23ffae7, 32'hc0d6cda3, 32'hc232c2cb, 32'hc2b81cbe};
test_label[2659] = '{32'h428b0da6};
test_output[2659] = '{32'h80000000};
/*############ DEBUG ############
test_input[21272:21279] = '{69.5266581757, -90.3409280116, -86.8281708636, -10.4742279786, -47.9950217544, -6.71260199812, -44.6902273355, -92.05613771};
test_label[2659] = '{69.5266581757};
test_output[2659] = '{-0.0};
############ END DEBUG ############*/
test_input[21280:21287] = '{32'h41853208, 32'h429d3ad4, 32'hc2ac2ecf, 32'hc101a828, 32'h42821065, 32'hc2c624b5, 32'hc288b8d5, 32'hc20df1df};
test_label[2660] = '{32'h41853208};
test_output[2660] = '{32'h4277dca4};
/*############ DEBUG ############
test_input[21280:21287] = '{16.6494301698, 78.6148967447, -86.091423596, -8.10355351606, 65.0320236831, -99.071696565, -68.3610004311, -35.4862038294};
test_label[2660] = '{16.6494301698};
test_output[2660] = '{61.9654678368};
############ END DEBUG ############*/
test_input[21288:21295] = '{32'h42089946, 32'h41c26998, 32'h42ada0ff, 32'hc0fc5f18, 32'h4146c249, 32'h41a4624c, 32'hc0e48f1b, 32'h428e2212};
test_label[2661] = '{32'h41c26998};
test_output[2661] = '{32'h427a0d33};
/*############ DEBUG ############
test_input[21288:21295] = '{34.1496819418, 24.3015595387, 86.8144485833, -7.88660827777, 12.4224324272, 20.5479971794, -7.14246873005, 71.066541889};
test_label[2661] = '{24.3015595387};
test_output[2661] = '{62.5128891894};
############ END DEBUG ############*/
test_input[21296:21303] = '{32'hc1940162, 32'hc1b852cd, 32'hc25c0cce, 32'hc13b918e, 32'h42bbf125, 32'h427d6087, 32'hc28afa0b, 32'hc2bcde70};
test_label[2662] = '{32'hc25c0cce};
test_output[2662] = '{32'h4314fbc6};
/*############ DEBUG ############
test_input[21296:21303] = '{-18.5006751646, -23.0404305987, -55.012506166, -11.7230357261, 93.9709876492, 63.3442658413, -69.4883684254, -94.4344447458};
test_label[2662] = '{-55.012506166};
test_output[2662] = '{148.983493815};
############ END DEBUG ############*/
test_input[21304:21311] = '{32'hc1e956bf, 32'hc2c4e3a5, 32'hc24fdbcb, 32'hc2a1c30a, 32'hc20e7595, 32'h3e74b51b, 32'hc1c3f9ef, 32'h423500c3};
test_label[2663] = '{32'hc20e7595};
test_output[2663] = '{32'h42a1bb2c};
/*############ DEBUG ############
test_input[21304:21311] = '{-29.1673569557, -98.4446167986, -51.9646423078, -80.8809387451, -35.6148261757, 0.238972116782, -24.4970380422, 45.2507423025};
test_label[2663] = '{-35.6148261757};
test_output[2663] = '{80.8655684783};
############ END DEBUG ############*/
test_input[21312:21319] = '{32'hc2a35375, 32'hc2a0ee22, 32'hc1e60c10, 32'h41e06ba4, 32'hc19e1396, 32'h4188decf, 32'hc13ad19d, 32'h42064585};
test_label[2664] = '{32'hc19e1396};
test_output[2664] = '{32'h4255536d};
/*############ DEBUG ############
test_input[21312:21319] = '{-81.6630032477, -80.4651032834, -28.7558897352, 28.0525590513, -19.7595634909, 17.1087925271, -11.676175388, 33.5678916628};
test_label[2664] = '{-19.7595634909};
test_output[2664] = '{53.331471736};
############ END DEBUG ############*/
test_input[21320:21327] = '{32'h420577fd, 32'h4254c08c, 32'h40bab48b, 32'hc1a96418, 32'h41a56d14, 32'h429ecf85, 32'hc284a604, 32'h40ee100d};
test_label[2665] = '{32'h4254c08c};
test_output[2665] = '{32'h41d1bcfb};
/*############ DEBUG ############
test_input[21320:21327] = '{33.3671752073, 53.1880351842, 5.83453900919, -21.1738744318, 20.6782602504, 79.4053103306, -66.3242482407, 7.43945923464};
test_label[2665] = '{53.1880351842};
test_output[2665] = '{26.2172751464};
############ END DEBUG ############*/
test_input[21328:21335] = '{32'h42a36840, 32'h3ee91fef, 32'hc28c6803, 32'h41743037, 32'h4291f263, 32'h42a62224, 32'hc226a0a0, 32'hc2be2d50};
test_label[2666] = '{32'h42a62224};
test_output[2666] = '{32'h3e695536};
/*############ DEBUG ############
test_input[21328:21335] = '{81.7036099073, 0.455321752703, -70.2031502069, 15.2617714857, 72.9734120638, 83.0666828244, -41.6568621666, -95.0885044136};
test_label[2666] = '{83.0666828244};
test_output[2666] = '{0.227864109637};
############ END DEBUG ############*/
test_input[21336:21343] = '{32'h414b13ae, 32'h425acaff, 32'h42a6abd5, 32'hc23bfe51, 32'h42a7936c, 32'hc23bac2c, 32'h42a722fb, 32'hc2b1cf4c};
test_label[2667] = '{32'h414b13ae};
test_output[2667] = '{32'h428ff973};
/*############ DEBUG ############
test_input[21336:21343] = '{12.6923043877, 54.6982398114, 83.3356079415, -46.998355253, 83.7879310094, -46.9181382625, 83.5683238976, -88.9048796207};
test_label[2667] = '{12.6923043877};
test_output[2667] = '{71.9872076795};
############ END DEBUG ############*/
test_input[21344:21351] = '{32'hc20e7308, 32'hc2b9ef78, 32'hc27baabd, 32'hc2b8bce4, 32'h427137fd, 32'h4285cf7b, 32'h402b77cc, 32'hc2a67e36};
test_label[2668] = '{32'h4285cf7b};
test_output[2668] = '{32'h3ab215f4};
/*############ DEBUG ############
test_input[21344:21351] = '{-35.6123363405, -92.9677142618, -62.9167356273, -92.36892498, 60.3046748242, 66.9052322909, 2.67918684093, -83.2465086086};
test_label[2668] = '{66.9052322909};
test_output[2668] = '{0.00135868645636};
############ END DEBUG ############*/
test_input[21352:21359] = '{32'hc1037fa5, 32'h420b9c1b, 32'h41322132, 32'hc2646252, 32'h422b5295, 32'h421876fb, 32'h4287f674, 32'hc255053e};
test_label[2669] = '{32'h4287f674};
test_output[2669] = '{32'h2d541880};
/*############ DEBUG ############
test_input[21352:21359] = '{-8.21866343968, 34.9024465052, 11.1331043417, -57.0960144755, 42.8306463058, 38.116192984, 67.9813555597, -53.2551184687};
test_label[2669] = '{67.9813555597};
test_output[2669] = '{1.20562448914e-11};
############ END DEBUG ############*/
test_input[21360:21367] = '{32'h42ae0469, 32'hc208781a, 32'hc2b9cd4d, 32'h41b41dd4, 32'hc253353d, 32'hc2a98c69, 32'h42398d39, 32'h424c96d0};
test_label[2670] = '{32'hc253353d};
test_output[2670] = '{32'h430bcf84};
/*############ DEBUG ############
test_input[21360:21367] = '{87.0086157639, -34.1172868999, -92.9009806165, 22.5145636134, -52.8019910492, -84.7742422397, 46.3879136907, 51.1472786297};
test_label[2670] = '{-52.8019910492};
test_output[2670] = '{139.810606813};
############ END DEBUG ############*/
test_input[21368:21375] = '{32'h3d8ebc81, 32'h42047b7b, 32'hbd8035b3, 32'h422f0442, 32'hc1d07e24, 32'hc2a45613, 32'h4279ea50, 32'hc25a85a8};
test_label[2671] = '{32'h42047b7b};
test_output[2671] = '{32'h41eaddaa};
/*############ DEBUG ############
test_input[21368:21375] = '{0.0696954769245, 33.1205878807, -0.0626024262936, 43.7541574325, -26.0615912285, -82.1681133445, 62.4788222014, -54.630522457};
test_label[2671] = '{33.1205878807};
test_output[2671] = '{29.358234328};
############ END DEBUG ############*/
test_input[21376:21383] = '{32'h4298cb58, 32'h42c1ffd8, 32'h424247ef, 32'h41cd4003, 32'hc28db763, 32'hc25f3093, 32'hc2932ace, 32'hc28ed1d6};
test_label[2672] = '{32'hc2932ace};
test_output[2672] = '{32'h432a9553};
/*############ DEBUG ############
test_input[21376:21383] = '{76.3971558774, 96.9996975438, 48.5702478905, 25.6562552585, -70.8581805566, -55.7974353536, -73.5836010938, -71.40983936};
test_label[2672] = '{-73.5836010938};
test_output[2672] = '{170.583298639};
############ END DEBUG ############*/
test_input[21384:21391] = '{32'h42c30d56, 32'h4250eacd, 32'h42bf74c4, 32'hc27f1247, 32'h429f5022, 32'h42362a12, 32'h42a5850f, 32'hc229c391};
test_label[2673] = '{32'hc27f1247};
test_output[2673] = '{32'h43217279};
/*############ DEBUG ############
test_input[21384:21391] = '{97.5260495787, 52.2292972281, 95.7280588523, -63.767849179, 79.656505682, 45.5410851563, 82.759880103, -42.4409845866};
test_label[2673] = '{-63.767849179};
test_output[2673] = '{161.447161978};
############ END DEBUG ############*/
test_input[21392:21399] = '{32'h4189168d, 32'hc1dd9b7f, 32'h41332d1c, 32'hc221fffb, 32'h4197c901, 32'hc1e5933c, 32'hc2a55759, 32'h421842ec};
test_label[2674] = '{32'hc1dd9b7f};
test_output[2674] = '{32'h42838855};
/*############ DEBUG ############
test_input[21392:21399] = '{17.1360118731, -27.7009255341, 11.1985133726, -40.4999810777, 18.9731458753, -28.6968924154, -82.6706026387, 38.0653515986};
test_label[2674] = '{-27.7009255341};
test_output[2674] = '{65.7662771387};
############ END DEBUG ############*/
test_input[21400:21407] = '{32'h4210e8fd, 32'h420e29d1, 32'hc29e93e9, 32'h429782cb, 32'hc27ee33b, 32'hc2c43ef1, 32'hc2c3c14c, 32'hc2c7cb13};
test_label[2675] = '{32'hc2c3c14c};
test_output[2675] = '{32'h432da20c};
/*############ DEBUG ############
test_input[21400:21407] = '{36.2275291205, 35.5408374031, -79.2888871542, 75.7554584816, -63.7219033877, -98.1229330315, -97.8775306866, -99.8966301448};
test_label[2675] = '{-97.8775306866};
test_output[2675] = '{173.632989168};
############ END DEBUG ############*/
test_input[21408:21415] = '{32'h42b51714, 32'h41c2bfcc, 32'h41f88053, 32'hc2a0fad9, 32'h3fb8a6f3, 32'hc1aa998b, 32'h41c31c8a, 32'h3f3b02b0};
test_label[2676] = '{32'hc2a0fad9};
test_output[2676] = '{32'h432b08f7};
/*############ DEBUG ############
test_input[21408:21415] = '{90.5450730904, 24.3436515418, 31.0626584724, -80.489939229, 1.44259483539, -21.3249724296, 24.3889354022, 0.730509740967};
test_label[2676] = '{-80.489939229};
test_output[2676] = '{171.035012319};
############ END DEBUG ############*/
test_input[21416:21423] = '{32'hc2868735, 32'hc28cdf65, 32'hc22e01e9, 32'hc1749c60, 32'h42711dc8, 32'h423a05ec, 32'h425ae4fd, 32'h42be1f95};
test_label[2677] = '{32'hc2868735};
test_output[2677] = '{32'h43225365};
/*############ DEBUG ############
test_input[21416:21423] = '{-67.2640770045, -70.4363146895, -43.5018666606, -15.2881778685, 60.2790848642, 46.505783283, 54.7236198879, 95.0616871684};
test_label[2677] = '{-67.2640770045};
test_output[2677] = '{162.325764173};
############ END DEBUG ############*/
test_input[21424:21431] = '{32'h4269c697, 32'h42ab107a, 32'h41aa1852, 32'hc14a74c8, 32'h41f1b2cd, 32'hc271eb71, 32'hc250346c, 32'h41bd0c0c};
test_label[2678] = '{32'hc271eb71};
test_output[2678] = '{32'h43120319};
/*############ DEBUG ############
test_input[21424:21431] = '{58.4439356802, 85.5321772975, 21.2618751578, -12.6535110922, 30.2123045579, -60.4799246382, -52.0511949516, 23.6308813646};
test_label[2678] = '{-60.4799246382};
test_output[2678] = '{146.012101936};
############ END DEBUG ############*/
test_input[21432:21439] = '{32'h42ac503d, 32'h4244af47, 32'hc28652a9, 32'hc23ea664, 32'h421efce0, 32'h4238dbec, 32'hc2565842, 32'h421f0be6};
test_label[2679] = '{32'hc28652a9};
test_output[2679] = '{32'h43195173};
/*############ DEBUG ############
test_input[21432:21439] = '{86.1567125667, 49.1711675857, -67.1614436177, -47.6624908405, 39.7469471662, 46.2147660661, -53.5861911471, 39.7616201518};
test_label[2679] = '{-67.1614436177};
test_output[2679] = '{153.318156184};
############ END DEBUG ############*/
test_input[21440:21447] = '{32'h42537e8d, 32'h42983dfc, 32'hc28f11de, 32'h4253ce10, 32'h4210ad4a, 32'hc2b78310, 32'h42a8266f, 32'hc2abdee5};
test_label[2680] = '{32'h4210ad4a};
test_output[2680] = '{32'h423f9fef};
/*############ DEBUG ############
test_input[21440:21447] = '{52.8735856282, 76.1210605757, -71.5348953893, 52.9512345014, 36.1692285542, -91.755978484, 84.0750626172, -85.935339538};
test_label[2680] = '{36.1692285542};
test_output[2680] = '{47.9061852549};
############ END DEBUG ############*/
test_input[21448:21455] = '{32'h416cbcb6, 32'h422e7734, 32'hc2b1eecb, 32'hc25a85ae, 32'h4217d461, 32'h421974ca, 32'hc23db9c2, 32'h4266c0f2};
test_label[2681] = '{32'h4266c0f2};
test_output[2681] = '{32'h35518377};
/*############ DEBUG ############
test_input[21448:21455] = '{14.7960720461, 43.616407863, -88.9663935238, -54.6305476786, 37.9573994453, 38.3640536569, -47.4314052395, 57.6884235434};
test_label[2681] = '{57.6884235434};
test_output[2681] = '{7.80498726149e-07};
############ END DEBUG ############*/
test_input[21456:21463] = '{32'h4158568d, 32'hc1d548ea, 32'hc29b063d, 32'h4140ff6e, 32'hc2744764, 32'hc28353da, 32'hc11f5dab, 32'h4281a8e9};
test_label[2682] = '{32'h4281a8e9};
test_output[2682] = '{32'h80000000};
/*############ DEBUG ############
test_input[21456:21463] = '{13.521130898, -26.6606017292, -77.5121811048, 12.0623609549, -61.0697182109, -65.6637757506, -9.9603682423, 64.8299001594};
test_label[2682] = '{64.8299001594};
test_output[2682] = '{-0.0};
############ END DEBUG ############*/
test_input[21464:21471] = '{32'hc28ba7eb, 32'hc24df354, 32'h42b8a3ad, 32'h429a4165, 32'hc2551eed, 32'h421503a4, 32'hc2955e27, 32'h42418479};
test_label[2683] = '{32'h421503a4};
test_output[2683] = '{32'h425c43b6};
/*############ DEBUG ############
test_input[21464:21471] = '{-69.8279647359, -51.4876236423, 92.3196780865, 77.1277254156, -53.280200683, 37.2535538414, -74.6838933552, 48.3793687996};
test_label[2683] = '{37.2535538414};
test_output[2683] = '{55.0661244976};
############ END DEBUG ############*/
test_input[21472:21479] = '{32'h42c4a7c6, 32'h429d10c9, 32'hc1e3955b, 32'hc2ba466a, 32'hc2c0d6ba, 32'hc29beb62, 32'h42c0ce3c, 32'hc18e0631};
test_label[2684] = '{32'h42c0ce3c};
test_output[2684] = '{32'h4003e882};
/*############ DEBUG ############
test_input[21472:21479] = '{98.3276822928, 78.5327828068, -28.4479274149, -93.1375288269, -96.4193904586, -77.9597324221, 96.4028005044, -17.7530236325};
test_label[2684] = '{96.4028005044};
test_output[2684] = '{2.06106603812};
############ END DEBUG ############*/
test_input[21480:21487] = '{32'hc04419f9, 32'h42bd9a50, 32'hc1120381, 32'hc0c6fe14, 32'hc1635c68, 32'h41cd47c4, 32'h423dc176, 32'hc2c1e3d6};
test_label[2685] = '{32'hc1635c68};
test_output[2685] = '{32'h42da05dd};
/*############ DEBUG ############
test_input[21480:21487] = '{-3.06408529352, 94.8013899015, -9.12585579873, -6.2185155366, -14.2100602445, 25.6600424792, 47.4389275954, -96.9449907739};
test_label[2685] = '{-14.2100602445};
test_output[2685] = '{109.011450146};
############ END DEBUG ############*/
test_input[21488:21495] = '{32'hc25b8722, 32'h40687197, 32'hbfb9c50d, 32'h41ea6dfa, 32'hc0e368f3, 32'h41ae9357, 32'h42100fb2, 32'h42a58d57};
test_label[2686] = '{32'h41ae9357};
test_output[2686] = '{32'h4273d103};
/*############ DEBUG ############
test_input[21488:21495] = '{-54.8819663033, 3.63193309134, -1.45132607107, 29.3036999821, -7.10656134278, 21.8219427414, 36.0153258386, 82.7760575713};
test_label[2686] = '{21.8219427414};
test_output[2686] = '{60.9541148299};
############ END DEBUG ############*/
test_input[21496:21503] = '{32'hc2a46edd, 32'hc16e1889, 32'hc28de924, 32'hc27ebc09, 32'h42033468, 32'h41844569, 32'hc18fed4d, 32'h41f356d1};
test_label[2687] = '{32'h42033468};
test_output[2687] = '{32'h3db49f7f};
/*############ DEBUG ############
test_input[21496:21503] = '{-82.2165315276, -14.8809900564, -70.9553544725, -63.683629833, 32.8011773128, 16.5338922977, -17.9908686183, 30.4173910487};
test_label[2687] = '{32.8011773128};
test_output[2687] = '{0.0881948395891};
############ END DEBUG ############*/
test_input[21504:21511] = '{32'hc2049c14, 32'hc2a52ea0, 32'h417c5c51, 32'h425af079, 32'hc2ab4519, 32'hc10ad0af, 32'hc1aa870f, 32'hc29b384d};
test_label[2688] = '{32'hc2ab4519};
test_output[2688] = '{32'h430c5eab};
/*############ DEBUG ############
test_input[21504:21511] = '{-33.15242157, -82.5910654432, 15.7725381945, 54.7348360847, -85.6349564525, -8.67594809165, -21.3159460232, -77.6099589892};
test_label[2688] = '{-85.6349564525};
test_output[2688] = '{140.369792537};
############ END DEBUG ############*/
test_input[21512:21519] = '{32'h421d31bc, 32'hc21e153e, 32'h429f75a2, 32'hc25a79ed, 32'hc220cb6b, 32'h413d5b14, 32'h42bdb302, 32'hc27f298a};
test_label[2689] = '{32'h413d5b14};
test_output[2689] = '{32'h42a607a0};
/*############ DEBUG ############
test_input[21512:21519] = '{39.2985696572, -39.520745263, 79.729748206, -54.6190700011, -40.1986519212, 11.8347356917, 94.8496262804, -63.7905646034};
test_label[2689] = '{11.8347356917};
test_output[2689] = '{83.0148908601};
############ END DEBUG ############*/
test_input[21520:21527] = '{32'h403ccce5, 32'hc2761256, 32'hbfdfdb85, 32'h40ac992b, 32'h4295989b, 32'h42c6e343, 32'h412e4b4f, 32'hc1a7e445};
test_label[2690] = '{32'hc2761256};
test_output[2690] = '{32'h4320f637};
/*############ DEBUG ############
test_input[21520:21527] = '{2.95000578601, -61.5179058052, -1.74888668919, 5.39369733008, 74.7980540105, 99.4438721516, 10.8933858706, -20.9864592286};
test_label[2690] = '{-61.5179058052};
test_output[2690] = '{160.961777957};
############ END DEBUG ############*/
test_input[21528:21535] = '{32'h41aff391, 32'h42a22651, 32'h420c1b18, 32'hc28a1bc6, 32'h428988ba, 32'h425ed27c, 32'h4103e601, 32'h4283e0f8};
test_label[2691] = '{32'h4103e601};
test_output[2691] = '{32'h4291a992};
/*############ DEBUG ############
test_input[21528:21535] = '{21.9939291969, 81.0748374384, 35.0264570719, -69.0542458299, 68.7670466552, 55.7055501201, 8.24365343776, 65.9393919471};
test_label[2691] = '{8.24365343776};
test_output[2691] = '{72.8311887843};
############ END DEBUG ############*/
test_input[21536:21543] = '{32'hc21760e4, 32'hc1520be3, 32'hc233f11b, 32'h415908aa, 32'hc2a8f766, 32'hc1d1d102, 32'hc219df18, 32'hc285fdbc};
test_label[2692] = '{32'hc1d1d102};
test_output[2692] = '{32'h421f2aac};
/*############ DEBUG ############
test_input[21536:21543] = '{-37.8446206869, -13.1279022484, -44.9854549941, 13.564615524, -84.4832008981, -26.2270545026, -38.4678637754, -66.9955752211};
test_label[2692] = '{-26.2270545026};
test_output[2692] = '{39.7916700266};
############ END DEBUG ############*/
test_input[21544:21551] = '{32'hc2c2a6a5, 32'h42286294, 32'hc226676d, 32'h40ab7320, 32'hc1f6b87f, 32'h4289d37c, 32'hc24853e3, 32'hbec31a1c};
test_label[2693] = '{32'hc1f6b87f};
test_output[2693] = '{32'h42c7819c};
/*############ DEBUG ############
test_input[21544:21551] = '{-97.32547478, 42.096267721, -41.600999948, 5.35780329638, -30.8400850413, 68.9130590089, -50.0819206273, -0.381058578099};
test_label[2693] = '{-30.8400850413};
test_output[2693] = '{99.7531440503};
############ END DEBUG ############*/
test_input[21552:21559] = '{32'h42146552, 32'hc2653647, 32'hc2b92901, 32'h42a490de, 32'h41aee728, 32'h41c2a4d4, 32'hc1b534b5, 32'hc28914da};
test_label[2694] = '{32'hc1b534b5};
test_output[2694] = '{32'h42d1de0b};
/*############ DEBUG ############
test_input[21552:21559] = '{37.0989466477, -57.3030054564, -92.5800860499, 82.2829456614, 21.8628690927, 24.3304823835, -22.6507353904, -68.5407233327};
test_label[2694] = '{-22.6507353904};
test_output[2694] = '{104.933681052};
############ END DEBUG ############*/
test_input[21560:21567] = '{32'hc2a9ef3e, 32'h42a69051, 32'h42a77994, 32'hc2533b2b, 32'h4265d71a, 32'hc217e098, 32'h42b15f0a, 32'hc1124334};
test_label[2695] = '{32'hc1124334};
test_output[2695] = '{32'h42c3ad58};
/*############ DEBUG ############
test_input[21560:21567] = '{-84.9672692325, 83.2818671245, 83.7374551278, -52.8077824258, 57.4600597938, -37.9693280875, 88.6856255201, -9.14140726436};
test_label[2695] = '{-9.14140726436};
test_output[2695] = '{97.8385620842};
############ END DEBUG ############*/
test_input[21568:21575] = '{32'h421f9c85, 32'h42adfe9d, 32'h4274ceaf, 32'hc2397434, 32'hc2354e44, 32'hc098afad, 32'hc14014c5, 32'hc245fa5c};
test_label[2696] = '{32'h42adfe9d};
test_output[2696] = '{32'h2cdc8f00};
/*############ DEBUG ############
test_input[21568:21575] = '{39.9028520344, 86.9972949169, 61.2018407582, -46.3634813824, -45.326429569, -4.77144480769, -12.005070306, -49.4944926679};
test_label[2696] = '{86.9972949169};
test_output[2696] = '{6.26865226396e-12};
############ END DEBUG ############*/
test_input[21576:21583] = '{32'hc2538354, 32'hc2add70e, 32'hc2c67a6a, 32'hc2a9d1bb, 32'h4201368f, 32'h42acd2e3, 32'hc21e021d, 32'hc2347c73};
test_label[2697] = '{32'h42acd2e3};
test_output[2697] = '{32'h80000000};
/*############ DEBUG ############
test_input[21576:21583] = '{-52.8782513615, -86.9200273282, -99.2390891425, -84.9096304108, 32.3032803677, 86.4118870294, -39.5020655117, -45.1215334882};
test_label[2697] = '{86.4118870294};
test_output[2697] = '{-0.0};
############ END DEBUG ############*/
test_input[21584:21591] = '{32'h42845dfe, 32'hc0c895eb, 32'hc2016ff7, 32'hc189eee7, 32'h420651a9, 32'h41cd3fb6, 32'h40ab72e5, 32'hc26565ae};
test_label[2698] = '{32'h40ab72e5};
test_output[2698] = '{32'h42734da0};
/*############ DEBUG ############
test_input[21584:21591] = '{66.1835809243, -6.26830061357, -32.3593403369, -17.2416510231, 33.5797472099, 25.6561087777, 5.35777533735, -57.3492951614};
test_label[2698] = '{5.35777533735};
test_output[2698] = '{60.825805587};
############ END DEBUG ############*/
test_input[21592:21599] = '{32'h428e8ac0, 32'h41efd87d, 32'h4291ac36, 32'h42b00bd6, 32'hc1f7f032, 32'hc1b07c7e, 32'h42ad15fe, 32'hc1f06b25};
test_label[2699] = '{32'h42ad15fe};
test_output[2699] = '{32'h3fd7b55c};
/*############ DEBUG ############
test_input[21592:21599] = '{71.2709978496, 29.9807079462, 72.8363493256, 88.0231143228, -30.9922819713, -22.0607862574, 86.5429545113, -30.0523165391};
test_label[2699] = '{86.5429545113};
test_output[2699] = '{1.68522217416};
############ END DEBUG ############*/
test_input[21600:21607] = '{32'hc2bc85c3, 32'h4171f29a, 32'h429ec2a1, 32'h42c675ab, 32'hc28d706c, 32'h424ad89d, 32'h420086b3, 32'hc2967b2c};
test_label[2700] = '{32'h4171f29a};
test_output[2700] = '{32'h42a83758};
/*############ DEBUG ############
test_input[21600:21607] = '{-94.2612521668, 15.1217287442, 79.3801313941, 99.2298192231, -70.7195711357, 50.7115362303, 32.1315433682, -75.2405695761};
test_label[2700] = '{15.1217287442};
test_output[2700] = '{84.1080904813};
############ END DEBUG ############*/
test_input[21608:21615] = '{32'hc2ae3757, 32'h4119ea66, 32'h42a365a0, 32'hc27d2cc5, 32'hc2008f77, 32'hc11bd632, 32'h3e9ab783, 32'hc2bee7ea};
test_label[2701] = '{32'hc2008f77};
test_output[2701] = '{32'h42e3ad5c};
/*############ DEBUG ############
test_input[21608:21615] = '{-87.1080825504, 9.61972652101, 81.6984877019, -63.2937210142, -32.1401016395, -9.73979367427, 0.302181328481, -95.4529533732};
test_label[2701] = '{-32.1401016395};
test_output[2701] = '{113.838589341};
############ END DEBUG ############*/
test_input[21616:21623] = '{32'hc191454a, 32'hc2ae8dbb, 32'hc247cbde, 32'hc2160fa1, 32'hc2449cb6, 32'h41627192, 32'hc2471109, 32'h42c09b2f};
test_label[2702] = '{32'hc2160fa1};
test_output[2702] = '{32'h4305d180};
/*############ DEBUG ############
test_input[21616:21623] = '{-18.1588327482, -87.276815127, -49.9490896647, -37.5152636255, -49.1530394337, 14.1527275676, -49.7666362642, 96.3030961243};
test_label[2702] = '{-37.5152636255};
test_output[2702] = '{133.81835975};
############ END DEBUG ############*/
test_input[21624:21631] = '{32'h428046da, 32'hc294dc04, 32'h4297055c, 32'h4268d328, 32'hc2753727, 32'hc2555c2f, 32'h42acb130, 32'hc1c44dee};
test_label[2703] = '{32'h4268d328};
test_output[2703] = '{32'h41e11e7b};
/*############ DEBUG ############
test_input[21624:21631] = '{64.1383797343, -74.4297203643, 75.510466352, 58.2062087349, -61.303860568, -53.3400240549, 86.3460711849, -24.5380516251};
test_label[2703] = '{58.2062087349};
test_output[2703] = '{28.139882136};
############ END DEBUG ############*/
test_input[21632:21639] = '{32'hc25e70ac, 32'h42186309, 32'hc2635487, 32'hc220012a, 32'hc1f18630, 32'h4250e2de, 32'hc28753ca, 32'hc2712daf};
test_label[2704] = '{32'hc220012a};
test_output[2704] = '{32'h42b87204};
/*############ DEBUG ############
test_input[21632:21639] = '{-55.6100293806, 38.0967158554, -56.8325447337, -40.0011363503, -30.1905220954, 52.221548983, -67.663653446, -60.2946136338};
test_label[2704] = '{-40.0011363503};
test_output[2704] = '{92.2226860673};
############ END DEBUG ############*/
test_input[21640:21647] = '{32'h41f861c7, 32'h4256395a, 32'h41ee70bf, 32'hc2936fa6, 32'hc296ac7c, 32'hc2ac8c9f, 32'h41d564fe, 32'h427c724e};
test_label[2705] = '{32'h427c724e};
test_output[2705] = '{32'h38947a3e};
/*############ DEBUG ############
test_input[21640:21647] = '{31.0477430354, 53.5560055576, 29.8050523147, -73.718064802, -75.3368838458, -86.2746469904, 26.6743124967, 63.1116274479};
test_label[2705] = '{63.1116274479};
test_output[2705] = '{7.07995941199e-05};
############ END DEBUG ############*/
test_input[21648:21655] = '{32'h41b24a8c, 32'hc07d1f8a, 32'hc2098a45, 32'h42348ed6, 32'hc195fbc8, 32'h4121abf6, 32'hc2a42b6c, 32'h42ac9060};
test_label[2706] = '{32'hc2a42b6c};
test_output[2706] = '{32'h43285de6};
/*############ DEBUG ############
test_input[21648:21655] = '{22.2864003986, -3.95504989733, -34.3850287607, 45.1394885887, -18.7479399179, 10.1044822859, -82.0848099539, 86.2819810951};
test_label[2706] = '{-82.0848099539};
test_output[2706] = '{168.366791049};
############ END DEBUG ############*/
test_input[21656:21663] = '{32'h411239a9, 32'h40c2c55d, 32'h42bcd0d3, 32'h420fbef2, 32'h41361498, 32'h4287e4eb, 32'hc27c68e3, 32'h42870384};
test_label[2707] = '{32'h420fbef2};
test_output[2707] = '{32'h4269e2b4};
/*############ DEBUG ############
test_input[21656:21663] = '{9.13907735785, 6.08659196957, 94.4078616704, 35.9364716765, 11.3800279572, 67.9471054873, -63.1024299816, 67.506868679};
test_label[2707] = '{35.9364716765};
test_output[2707] = '{58.4713899939};
############ END DEBUG ############*/
test_input[21664:21671] = '{32'hc2b49e85, 32'hc2b086c3, 32'hc2ba5dc6, 32'h42c65458, 32'hc291bd31, 32'h41975654, 32'h42818d7f, 32'hc2a97a33};
test_label[2708] = '{32'hc2b086c3};
test_output[2708] = '{32'h433b6d8d};
/*############ DEBUG ############
test_input[21664:21671] = '{-90.3096082631, -88.2632060039, -93.1831546155, 99.1647319067, -72.8695170359, 18.9171527543, 64.7763631184, -84.7386685408};
test_label[2708] = '{-88.2632060039};
test_output[2708] = '{187.427937911};
############ END DEBUG ############*/
test_input[21672:21679] = '{32'h41e4abe5, 32'hc156bebe, 32'hc2900227, 32'h40d476ef, 32'hc2887ca4, 32'hc2b2dc09, 32'hc2a16b9b, 32'h42b57eb4};
test_label[2709] = '{32'hc2b2dc09};
test_output[2709] = '{32'h43342d5e};
/*############ DEBUG ############
test_input[21672:21679] = '{28.5839324121, -13.4215683553, -72.0042029781, 6.63951812094, -68.2434389344, -89.4297536803, -80.7101648141, 90.7474669093};
test_label[2709] = '{-89.4297536803};
test_output[2709] = '{180.17722059};
############ END DEBUG ############*/
test_input[21680:21687] = '{32'h42c21ce6, 32'hc19fdd0c, 32'h420dd108, 32'h42672466, 32'hc1d5510a, 32'h4287fff3, 32'h429d534e, 32'hc26815b6};
test_label[2710] = '{32'hc26815b6};
test_output[2710] = '{32'h431b13e1};
/*############ DEBUG ############
test_input[21680:21687] = '{97.0564434527, -19.9829327444, 35.4541317654, 57.7855436656, -26.6645699494, 67.9999005976, 78.662707359, -58.0212030401};
test_label[2710] = '{-58.0212030401};
test_output[2710] = '{155.077646503};
############ END DEBUG ############*/
test_input[21688:21695] = '{32'h421c135d, 32'hc1cc0f0d, 32'hc2a7184b, 32'hc17ff7cd, 32'hc28172c2, 32'hc2bafae9, 32'hc28ee222, 32'h428c417a};
test_label[2711] = '{32'h421c135d};
test_output[2711] = '{32'h41f8df2c};
/*############ DEBUG ############
test_input[21688:21695] = '{39.0189100609, -25.5073487957, -83.5474479195, -15.9979980563, -64.7241386129, -93.4900594884, -71.4416629864, 70.1278805785};
test_label[2711] = '{39.0189100609};
test_output[2711] = '{31.1089705176};
############ END DEBUG ############*/
test_input[21696:21703] = '{32'h42c15099, 32'h422b247e, 32'h42351c7e, 32'h429a310e, 32'hc1c2ea2f, 32'hc2a71130, 32'hc2813913, 32'hc292a1c0};
test_label[2712] = '{32'hc2a71130};
test_output[2712] = '{32'h433430e5};
/*############ DEBUG ############
test_input[21696:21703] = '{96.6574157301, 42.7856352176, 45.277824001, 77.0958134025, -24.3643483819, -83.5335710322, -64.6114766485, -73.3159199539};
test_label[2712] = '{-83.5335710322};
test_output[2712] = '{180.190986766};
############ END DEBUG ############*/
test_input[21704:21711] = '{32'hc2536754, 32'hc0dbec45, 32'h4190a455, 32'hc27cc8f6, 32'hc18bd8d0, 32'h42a5082b, 32'hc2489b8a, 32'hc28c1cb5};
test_label[2713] = '{32'hc28c1cb5};
test_output[2713] = '{32'h43189270};
/*############ DEBUG ############
test_input[21704:21711] = '{-52.8509045361, -6.872591493, 18.0802408483, -63.1962515607, -17.4808658897, 82.5159526577, -50.1518926551, -70.056066188};
test_label[2713] = '{-70.056066188};
test_output[2713] = '{152.572018846};
############ END DEBUG ############*/
test_input[21712:21719] = '{32'hc1c74bd3, 32'h419107a8, 32'h42206047, 32'h42958e5d, 32'hc161ef86, 32'h4015dc8c, 32'h41b12ada, 32'hc29076cc};
test_label[2714] = '{32'h4015dc8c};
test_output[2714] = '{32'h4290df78};
/*############ DEBUG ############
test_input[21712:21719] = '{-24.9120231264, 18.1287376354, 40.0940213152, 74.7780514242, -14.1209776824, 2.34158617031, 22.1459242542, -72.2320264974};
test_label[2714] = '{2.34158617031};
test_output[2714] = '{72.4364652539};
############ END DEBUG ############*/
test_input[21720:21727] = '{32'h42a21839, 32'h40c4d12c, 32'hc0b63e54, 32'hc22ee249, 32'h42bb7c86, 32'hc20b6409, 32'hc1f90378, 32'h42c263f4};
test_label[2715] = '{32'hc20b6409};
test_output[2715] = '{32'h430412f8};
/*############ DEBUG ############
test_input[21720:21727] = '{81.0473093778, 6.15053360092, -5.69510833989, -43.7209809698, 93.7432067639, -34.8476897367, -31.1266938425, 97.1952171646};
test_label[2715] = '{-34.8476897367};
test_output[2715] = '{132.074097358};
############ END DEBUG ############*/
test_input[21728:21735] = '{32'h42bc8ae9, 32'hc0e3d9da, 32'h42c25cfc, 32'h4281a15f, 32'h409f6d7c, 32'hc20eebd7, 32'hc29ca2b9, 32'hc0a8a23e};
test_label[2716] = '{32'hc0e3d9da};
test_output[2716] = '{32'h42d0b5c0};
/*############ DEBUG ############
test_input[21728:21735] = '{94.2713106595, -7.12034336175, 97.1816093676, 64.8151749296, 4.9821146077, -35.7303122064, -78.3178155682, -5.26980509728};
test_label[2716] = '{-7.12034336175};
test_output[2716] = '{104.354981005};
############ END DEBUG ############*/
test_input[21736:21743] = '{32'hc2c5710f, 32'hc23fd932, 32'h4210de56, 32'h42361520, 32'h403cc865, 32'hc26d3f55, 32'h413d7319, 32'h42046074};
test_label[2717] = '{32'h42046074};
test_output[2717] = '{32'h4146d315};
/*############ DEBUG ############
test_input[21736:21743] = '{-98.7208196146, -47.9621064499, 36.2171239338, 45.5206307473, 2.9497310894, -59.3118469648, 11.8405996589, 33.0941919441};
test_label[2717] = '{33.0941919441};
test_output[2717] = '{12.426533914};
############ END DEBUG ############*/
test_input[21744:21751] = '{32'hc2351e78, 32'h42bb710f, 32'hc20b546b, 32'h427ef425, 32'hc1763bcf, 32'hc25036e4, 32'hc2aab521, 32'h41a7a2be};
test_label[2718] = '{32'hc20b546b};
test_output[2718] = '{32'h43008da3};
/*############ DEBUG ############
test_input[21744:21751] = '{-45.2797527542, 93.7208208389, -34.8324405158, 63.7384228034, -15.3896019053, -52.0536045747, -85.3537646111, 20.9544638056};
test_label[2718] = '{-34.8324405158};
test_output[2718] = '{128.553261355};
############ END DEBUG ############*/
test_input[21752:21759] = '{32'h428c1730, 32'h424472cc, 32'hc28eb492, 32'hc19e1808, 32'hc0b7a5b6, 32'h42bfb07f, 32'h42c4ea6f, 32'h42a78e5b};
test_label[2719] = '{32'h428c1730};
test_output[2719] = '{32'h41e3dddf};
/*############ DEBUG ############
test_input[21752:21759] = '{70.0452850008, 49.1121044175, -71.352673594, -19.7617346233, -5.73897860978, 95.8447182297, 98.4578792913, 83.7780374053};
test_label[2719] = '{70.0452850008};
test_output[2719] = '{28.4833349928};
############ END DEBUG ############*/
test_input[21760:21767] = '{32'hc216d1e0, 32'h42bccf38, 32'hc29f38ed, 32'hc15a5372, 32'h4243c6b7, 32'hc2c02c9b, 32'hc2b2339d, 32'h41aad2c2};
test_label[2720] = '{32'hc216d1e0};
test_output[2720] = '{32'h43041c14};
/*############ DEBUG ############
test_input[21760:21767] = '{-37.7049572104, 94.4047254355, -79.6111818919, -13.6453721145, 48.9440580756, -96.0871233786, -89.1008095132, 21.3529082189};
test_label[2720] = '{-37.7049572104};
test_output[2720] = '{132.109682646};
############ END DEBUG ############*/
test_input[21768:21775] = '{32'h42c5a0bb, 32'hc273d43d, 32'h4289de84, 32'h408cf96d, 32'h429fd158, 32'h426f04b2, 32'hc1901bd0, 32'h3fbc33f6};
test_label[2721] = '{32'h426f04b2};
test_output[2721] = '{32'h421c3cc3};
/*############ DEBUG ############
test_input[21768:21775] = '{98.8139241554, -60.9572656703, 68.9346039318, 4.40544749274, 79.908877377, 59.7545866113, -18.0135807133, 1.4703357263};
test_label[2721] = '{59.7545866113};
test_output[2721] = '{39.0593375503};
############ END DEBUG ############*/
test_input[21776:21783] = '{32'hc29dc068, 32'h41c81926, 32'h42bbed48, 32'hc22b9254, 32'hc276257b, 32'hc25c9743, 32'hc2a4af7e, 32'hc2ab75b3};
test_label[2722] = '{32'hc2ab75b3};
test_output[2722] = '{32'h4333b17e};
/*############ DEBUG ############
test_input[21776:21783] = '{-78.8757953015, 25.0122787922, 93.9634368739, -42.8928983999, -61.5366024974, -55.1477170346, -82.3427564275, -85.7298850175};
test_label[2722] = '{-85.7298850175};
test_output[2722] = '{179.693321891};
############ END DEBUG ############*/
test_input[21784:21791] = '{32'h41fedc5e, 32'h4248cc19, 32'h426c909e, 32'hc2c152a0, 32'h42a00d8a, 32'h411a6e60, 32'h42473edc, 32'hc246dc1d};
test_label[2723] = '{32'h426c909e};
test_output[2723] = '{32'h41a714ed};
/*############ DEBUG ############
test_input[21784:21791] = '{31.8576005684, 50.1993122741, 59.1412269643, -96.6613790213, 80.0264451285, 9.65194704073, 49.8113874481, -49.7149549308};
test_label[2723] = '{59.1412269643};
test_output[2723] = '{20.8852181651};
############ END DEBUG ############*/
test_input[21792:21799] = '{32'h413699f6, 32'h42918885, 32'h420c2ef3, 32'h42aa775d, 32'h42959ad4, 32'hc20331dc, 32'h4196d6f9, 32'hc08bd95e};
test_label[2724] = '{32'h42918885};
test_output[2724] = '{32'h414776e5};
/*############ DEBUG ############
test_input[21792:21799] = '{11.4125880011, 72.7666388949, 35.0458495261, 85.233132258, 74.8023989937, -32.7986898139, 18.8549664017, -4.37028394515};
test_label[2724] = '{72.7666388949};
test_output[2724] = '{12.4665267276};
############ END DEBUG ############*/
test_input[21800:21807] = '{32'h41cdfd77, 32'h42a541ca, 32'h42959a4e, 32'h424ab7c2, 32'hc169c9e8, 32'h4258216c, 32'hc21f6fa1, 32'h42b05e6a};
test_label[2725] = '{32'h41cdfd77};
test_output[2725] = '{32'h4279c20c};
/*############ DEBUG ############
test_input[21800:21807] = '{25.7487623099, 82.628491393, 74.8013739247, 50.679451904, -14.6117936023, 54.0326394756, -39.859012016, 88.1844024272};
test_label[2725] = '{25.7487623099};
test_output[2725] = '{62.4394987504};
############ END DEBUG ############*/
test_input[21808:21815] = '{32'h42725644, 32'h41e6b501, 32'h42553d36, 32'h42ab751b, 32'hc272d7f3, 32'hc2452ab4, 32'hc2b392db, 32'h422097b7};
test_label[2726] = '{32'hc2452ab4};
test_output[2726] = '{32'h4307053b};
/*############ DEBUG ############
test_input[21808:21815] = '{60.5842442149, 28.8383811201, 53.3097782032, 85.7287245132, -60.7108868971, -49.2917031469, -89.7868254272, 40.1481591472};
test_label[2726] = '{-49.2917031469};
test_output[2726] = '{135.02042766};
############ END DEBUG ############*/
test_input[21816:21823] = '{32'h3fc90366, 32'h42ada378, 32'h42b265ee, 32'h3f4fa8d2, 32'h409930ec, 32'hc2bba0a0, 32'h411616b8, 32'h42155825};
test_label[2727] = '{32'h42155825};
test_output[2727] = '{32'h424fce60};
/*############ DEBUG ############
test_input[21816:21823] = '{1.57041617962, 86.819274501, 89.1990836804, 0.811169758905, 4.78722214495, -93.8137190921, 9.38054652501, 37.3360775485};
test_label[2727] = '{37.3360775485};
test_output[2727] = '{51.9515372399};
############ END DEBUG ############*/
test_input[21824:21831] = '{32'hc29184b1, 32'hc209a869, 32'h414a06a7, 32'hc1938ade, 32'h4147f53b, 32'hc19c7e69, 32'hc253df52, 32'h41542655};
test_label[2728] = '{32'h41542655};
test_output[2728] = '{32'h3f312c71};
/*############ DEBUG ############
test_input[21824:21831] = '{-72.7591644755, -34.4144616982, 12.6266243174, -18.4428065036, 12.4973707571, -19.5617236608, -52.9680880196, 13.2593583713};
test_label[2728] = '{13.2593583713};
test_output[2728] = '{0.692084348373};
############ END DEBUG ############*/
test_input[21832:21839] = '{32'hc2b6c808, 32'h422613c1, 32'hc2a6aebc, 32'h41a54686, 32'hc2022134, 32'h42288c0a, 32'hc16365a9, 32'hc2b6850c};
test_label[2729] = '{32'h41a54686};
test_output[2729] = '{32'h41af44ec};
/*############ DEBUG ############
test_input[21832:21839] = '{-91.3906863495, 41.519291697, -83.3412745395, 20.6594359932, -32.5324236737, 42.1367551018, -14.2123191396, -91.2598583064};
test_label[2729] = '{20.6594359932};
test_output[2729] = '{21.9086538388};
############ END DEBUG ############*/
test_input[21840:21847] = '{32'h428ec350, 32'h4287fdd8, 32'hc1b7b2f0, 32'hbf6d3ea8, 32'hbf25ccb5, 32'hc2a3b031, 32'hc2c72661, 32'hc1588ddf};
test_label[2730] = '{32'h4287fdd8};
test_output[2730] = '{32'h405ad088};
/*############ DEBUG ############
test_input[21840:21847] = '{71.3814688927, 67.9957852144, -22.9623723273, -0.926737312626, -0.64765483284, -81.8441202518, -99.5749605067, -13.5346362128};
test_label[2730] = '{67.9957852144};
test_output[2730] = '{3.41897771797};
############ END DEBUG ############*/
test_input[21848:21855] = '{32'h422c17d1, 32'hc2a5b326, 32'h41f64de1, 32'h4283f179, 32'hc19abe6b, 32'hc01fbc09, 32'hc28d4bcf, 32'h4291514e};
test_label[2731] = '{32'hc01fbc09};
test_output[2731] = '{32'h42964fd2};
/*############ DEBUG ############
test_input[21848:21855] = '{43.0232573527, -82.8498974908, 30.7880264406, 65.9716277286, -19.3429783015, -2.4958516911, -70.6480660736, 72.6588014482};
test_label[2731] = '{-2.4958516911};
test_output[2731] = '{75.1558991643};
############ END DEBUG ############*/
test_input[21856:21863] = '{32'h42c23a88, 32'h4218a2aa, 32'h41ee8401, 32'h42b3134c, 32'h417761ee, 32'h428a1a09, 32'h4263e5a1, 32'hc27ebf3e};
test_label[2732] = '{32'h428a1a09};
test_output[2732] = '{32'h41e0830a};
/*############ DEBUG ############
test_input[21856:21863] = '{97.1143222095, 38.1588517441, 29.8144554099, 89.5376917421, 15.4614090866, 69.050850781, 56.974246191, -63.6867616522};
test_label[2732] = '{69.050850781};
test_output[2732] = '{28.0639835818};
############ END DEBUG ############*/
test_input[21864:21871] = '{32'hc1442aaf, 32'hc2c1a2cd, 32'hc2863eb7, 32'h42bb2db4, 32'h42b4abc1, 32'hc23755a2, 32'h41d48220, 32'hc1c90cf8};
test_label[2733] = '{32'h42b4abc1};
test_output[2733] = '{32'h4052ab5f};
/*############ DEBUG ############
test_input[21864:21871] = '{-12.2604205613, -96.8179715577, -67.1224926311, 93.5892634316, 90.3354532951, -45.8336266455, 26.5635374214, -25.1313323479};
test_label[2733] = '{90.3354532951};
test_output[2733] = '{3.29170954821};
############ END DEBUG ############*/
test_input[21872:21879] = '{32'h41b5344c, 32'h41670e5c, 32'hc2537449, 32'h420a637a, 32'hc2b4a58f, 32'hc1946406, 32'h40f0c483, 32'hc22b05c3};
test_label[2734] = '{32'hc2537449};
test_output[2734] = '{32'h42aeebe2};
/*############ DEBUG ############
test_input[21872:21879] = '{22.6505352628, 14.4410055552, -52.8635582792, 34.597144807, -90.3233568248, -18.5488402729, 7.52398826331, -42.7556258711};
test_label[2734] = '{-52.8635582792};
test_output[2734] = '{87.4607095691};
############ END DEBUG ############*/
test_input[21880:21887] = '{32'hc2ae5766, 32'h4132c938, 32'hc2399d4c, 32'hc1f7e282, 32'h415c0e3e, 32'h42b42f81, 32'hc2c11912, 32'h40becc38};
test_label[2735] = '{32'h415c0e3e};
test_output[2735] = '{32'h4298adb9};
/*############ DEBUG ############
test_input[21880:21887] = '{-87.1706970334, 11.1741260254, -46.4036098632, -30.9855990079, 13.7534771909, 90.0927802381, -96.5489650133, 5.96242894158};
test_label[2735] = '{13.7534771909};
test_output[2735] = '{76.3393030472};
############ END DEBUG ############*/
test_input[21888:21895] = '{32'h42331346, 32'hc2872bcb, 32'h4281fcf0, 32'h4217d3fc, 32'h41da7dc2, 32'h4293fd0c, 32'h427857ea, 32'hc1ef04dc};
test_label[2736] = '{32'h4217d3fc};
test_output[2736] = '{32'h4210263f};
/*############ DEBUG ############
test_input[21888:21895] = '{44.7688216454, -67.5855336872, 64.9940204849, 37.9570143336, 27.3114049416, 73.9942323874, 62.0858542943, -29.8773720933};
test_label[2736] = '{37.9570143336};
test_output[2736] = '{36.0373481628};
############ END DEBUG ############*/
test_input[21896:21903] = '{32'h4208b7c1, 32'h41a656da, 32'hc2b73500, 32'h420e125b, 32'h427ce953, 32'hc2053a7c, 32'hbf61dfb2, 32'hc26706ba};
test_label[2737] = '{32'h4208b7c1};
test_output[2737] = '{32'h41e86325};
/*############ DEBUG ############
test_input[21896:21903] = '{34.1794469994, 20.7924079097, -91.6035132608, 35.5179261757, 63.2278565505, -33.3071122364, -0.882319587103, -57.7565682275};
test_label[2737] = '{34.1794469994};
test_output[2737] = '{29.0484095511};
############ END DEBUG ############*/
test_input[21904:21911] = '{32'hc26744fe, 32'hc2343837, 32'h422d931c, 32'hc1ba16b9, 32'hc2b5a64f, 32'h424c690a, 32'hc17dfce3, 32'h41d3bc70};
test_label[2738] = '{32'hc1ba16b9};
test_output[2738] = '{32'h4294ba6e};
/*############ DEBUG ############
test_input[21904:21911] = '{-57.8173756551, -45.0548959159, 43.3936615751, -23.2610953084, -90.8248226541, 51.102577579, -15.8742396164, 26.4670114245};
test_label[2738] = '{-23.2610953084};
test_output[2738] = '{74.3641215945};
############ END DEBUG ############*/
test_input[21912:21919] = '{32'h420b67c6, 32'h425375be, 32'h425aee18, 32'h428c4162, 32'hc0a5bc97, 32'hc144be31, 32'h411b1427, 32'hc236976e};
test_label[2739] = '{32'hc236976e};
test_output[2739] = '{32'h42e78d18};
/*############ DEBUG ############
test_input[21912:21919] = '{34.8513403921, 52.8649844577, 54.7325135321, 70.1276975585, -5.17927137656, -12.296433384, 9.69241962728, -45.6478788661};
test_label[2739] = '{-45.6478788661};
test_output[2739] = '{115.775576662};
############ END DEBUG ############*/
test_input[21920:21927] = '{32'h42a41544, 32'h42b48d54, 32'h4263b6bd, 32'h424cc194, 32'hc154f9f4, 32'hc1470854, 32'h429db470, 32'h42beece6};
test_label[2740] = '{32'hc1470854};
test_output[2740] = '{32'h42d7d0cc};
/*############ DEBUG ############
test_input[21920:21927] = '{82.0415351846, 90.2760288976, 56.9284568319, 51.1890412363, -13.3110239134, -12.4395331848, 78.8524155091, 95.4626936813};
test_label[2740] = '{-12.4395331848};
test_output[2740] = '{107.907803454};
############ END DEBUG ############*/
test_input[21928:21935] = '{32'h42af4862, 32'hc1d8ad68, 32'h41531200, 32'h42928850, 32'h428f05f9, 32'h42a89f24, 32'hc246fec1, 32'h4252bbcd};
test_label[2741] = '{32'h41531200};
test_output[2741] = '{32'h4294f821};
/*############ DEBUG ############
test_input[21928:21935] = '{87.641374398, -27.0846713795, 13.1918945099, 73.2662315833, 71.5116666223, 84.3108223535, -49.748782026, 52.6833988305};
test_label[2741] = '{13.1918945099};
test_output[2741] = '{74.4846288821};
############ END DEBUG ############*/
test_input[21936:21943] = '{32'h4120b3d7, 32'h4152f1d2, 32'h40baaed1, 32'h40a6665a, 32'h425d4b93, 32'h4293cdd9, 32'hc213c658, 32'hc2233dc8};
test_label[2742] = '{32'h40baaed1};
test_output[2742] = '{32'h428822ec};
/*############ DEBUG ############
test_input[21936:21943] = '{10.0439057513, 13.1840379239, 5.83383986549, 5.19999422527, 55.3238020207, 73.902044053, -36.9436953081, -40.8103323572};
test_label[2742] = '{5.83383986549};
test_output[2742] = '{68.0682041961};
############ END DEBUG ############*/
test_input[21944:21951] = '{32'hc2869e31, 32'hc265abfc, 32'h41c0557a, 32'h42637e8c, 32'h42b2ce86, 32'hc2ac8600, 32'h4226a245, 32'hc1f87331};
test_label[2743] = '{32'h42b2ce86};
test_output[2743] = '{32'h28060000};
/*############ DEBUG ############
test_input[21944:21951] = '{-67.3089693291, -57.4179528277, 24.041735993, 56.8735800307, 89.4033686597, -86.2617180186, 41.6584680631, -31.0562458166};
test_label[2743] = '{89.4033686597};
test_output[2743] = '{7.43849426499e-15};
############ END DEBUG ############*/
test_input[21952:21959] = '{32'hc2be76ba, 32'hc1ff2372, 32'hc228d8bc, 32'hc2683ce0, 32'h412e6657, 32'hc14f404a, 32'hc296da02, 32'hc0370474};
test_label[2744] = '{32'hc2be76ba};
test_output[2744] = '{32'h42d44385};
/*############ DEBUG ############
test_input[21952:21959] = '{-95.2318865064, -31.8923076075, -42.2116538661, -58.0594491901, 10.8999855939, -12.9531960013, -75.4257936163, -2.85964679702};
test_label[2744] = '{-95.2318865064};
test_output[2744] = '{106.131873158};
############ END DEBUG ############*/
test_input[21960:21967] = '{32'h41a104d1, 32'hc2aced09, 32'hc2adec91, 32'hc28f7e74, 32'hc1d46705, 32'hc2092108, 32'hc2a8da2f, 32'hc28eac83};
test_label[2745] = '{32'h41a104d1};
test_output[2745] = '{32'h80000000};
/*############ DEBUG ############
test_input[21960:21967] = '{20.1273521025, -86.462959392, -86.9620436177, -71.7469778716, -26.5503018414, -34.2822589821, -84.426139955, -71.3369337667};
test_label[2745] = '{20.1273521025};
test_output[2745] = '{-0.0};
############ END DEBUG ############*/
test_input[21968:21975] = '{32'h4003358d, 32'h3c32a518, 32'hc13b43f2, 32'h42b8727d, 32'hc2b909ae, 32'hc21aa41e, 32'hc237e825, 32'hc229982e};
test_label[2746] = '{32'h42b8727d};
test_output[2746] = '{32'h80000000};
/*############ DEBUG ############
test_input[21968:21975] = '{2.05014358512, 0.0109036192222, -11.7040884843, 92.2236072426, -92.5189026363, -38.6602723444, -45.9767028141, -42.3986146005};
test_label[2746] = '{92.2236072426};
test_output[2746] = '{-0.0};
############ END DEBUG ############*/
test_input[21976:21983] = '{32'hc23ccd7a, 32'hc1cfaa2a, 32'hc2896a16, 32'h426cac7c, 32'h422c6b4e, 32'hc1b0b3ec, 32'h42a719d6, 32'h41aea00d};
test_label[2747] = '{32'h42a719d6};
test_output[2747] = '{32'h2de2a080};
/*############ DEBUG ############
test_input[21976:21983] = '{-47.2006597785, -25.9580883553, -68.7071980869, 59.1684407423, 43.104788411, -22.0878533848, 83.5504636056, 21.8281497973};
test_label[2747] = '{83.5504636056};
test_output[2747] = '{2.57645016436e-11};
############ END DEBUG ############*/
test_input[21984:21991] = '{32'hc1504553, 32'h42255837, 32'hc1a00faf, 32'h41f6cf9e, 32'hc2094a8f, 32'hc18fd1ce, 32'hc2993d60, 32'h42825857};
test_label[2748] = '{32'h42255837};
test_output[2748] = '{32'h41beb0ee};
/*############ DEBUG ############
test_input[21984:21991] = '{-13.0169247052, 41.3361468008, -20.0076572652, 30.8513762749, -34.3228121031, -17.977444125, -76.6198695174, 65.1725386369};
test_label[2748] = '{41.3361468008};
test_output[2748] = '{23.8363918362};
############ END DEBUG ############*/
test_input[21992:21999] = '{32'hc2896395, 32'hc2975e43, 32'hc2c506de, 32'h3eeb67f8, 32'hc29f53fc, 32'hc2ad695f, 32'hc28b8e32, 32'hc2a81708};
test_label[2749] = '{32'hc29f53fc};
test_output[2749] = '{32'h42a03f64};
/*############ DEBUG ############
test_input[21992:21999] = '{-68.6944986393, -75.6841019386, -98.5134132807, 0.459777596449, -79.6640317669, -86.7057998516, -69.777724731, -84.0449791988};
test_label[2749] = '{-79.6640317669};
test_output[2749] = '{80.1238093634};
############ END DEBUG ############*/
test_input[22000:22007] = '{32'h424bfb5c, 32'h4230e7ed, 32'h429efad1, 32'hc1c09e2d, 32'h4229eb16, 32'h42489140, 32'h4265fb51, 32'h418603a5};
test_label[2750] = '{32'h424bfb5c};
test_output[2750] = '{32'h41e3f48c};
/*############ DEBUG ############
test_input[22000:22007] = '{50.9954665037, 44.2264892008, 79.4898740348, -24.0772350095, 42.479577579, 50.1418464015, 57.4954259517, 16.7517804844};
test_label[2750] = '{50.9954665037};
test_output[2750] = '{28.4944075314};
############ END DEBUG ############*/
test_input[22008:22015] = '{32'hc29ef1b0, 32'hc284c13d, 32'h42bdf40f, 32'h422d04cd, 32'h42c00463, 32'h3facb50c, 32'hc1350bbd, 32'h4279edc0};
test_label[2751] = '{32'hc284c13d};
test_output[2751] = '{32'h4322b0d6};
/*############ DEBUG ############
test_input[22008:22015] = '{-79.4720449847, -66.3774149509, 94.9766733838, 43.2546884307, 96.0085704772, 1.34927513107, -11.3153661186, 62.4821777266};
test_label[2751] = '{-66.3774149509};
test_output[2751] = '{162.690768192};
############ END DEBUG ############*/
test_input[22016:22023] = '{32'h429a6980, 32'hc286a1f3, 32'hc2110748, 32'hc2885848, 32'h4289ac5c, 32'hc29a0735, 32'h40883cee, 32'hc22c7f42};
test_label[2752] = '{32'h40883cee};
test_output[2752] = '{32'h4291e5cf};
/*############ DEBUG ############
test_input[22016:22023] = '{77.2060513431, -67.3163084264, -36.2571108025, -68.1724220481, 68.8366388634, -77.0140761641, 4.25743770462, -43.1242744984};
test_label[2752] = '{4.25743770462};
test_output[2752] = '{72.9488454633};
############ END DEBUG ############*/
test_input[22024:22031] = '{32'h42b43c0b, 32'h41ef5526, 32'h422f657b, 32'hc2a43e37, 32'h40fa36ec, 32'hc10f1819, 32'hc1f8de2e, 32'hc24065ed};
test_label[2753] = '{32'h422f657b};
test_output[2753] = '{32'h4239129c};
/*############ DEBUG ############
test_input[22024:22031] = '{90.1172744035, 29.9165767661, 43.849102595, -82.1215164993, 7.81920425931, -8.94338301028, -31.1084856728, -48.0995371086};
test_label[2753] = '{43.849102595};
test_output[2753] = '{46.2681718085};
############ END DEBUG ############*/
test_input[22032:22039] = '{32'h41a9f1f5, 32'hc1f99157, 32'h42505116, 32'h42178b7a, 32'h427a4a6f, 32'hc27fb314, 32'hc1aa857c, 32'hc206e23d};
test_label[2754] = '{32'hc206e23d};
test_output[2754] = '{32'h42c0965a};
/*############ DEBUG ############
test_input[22032:22039] = '{21.2431439949, -31.1959667273, 52.0791869003, 37.8862084109, 62.5726884822, -63.9248811498, -21.3151774906, -33.7209364568};
test_label[2754] = '{-33.7209364568};
test_output[2754] = '{96.2936526547};
############ END DEBUG ############*/
test_input[22040:22047] = '{32'hc149364a, 32'hc1ed724e, 32'h42c4ba6d, 32'h42adc8bd, 32'h42c0b6f1, 32'hc13a4bc4, 32'hc233acf1, 32'h429c2151};
test_label[2755] = '{32'h42c0b6f1};
test_output[2755] = '{32'h400881fe};
/*############ DEBUG ############
test_input[22040:22047] = '{-12.5757537362, -29.6808124195, 98.364110372, 86.8920639536, 96.3573047515, -11.6434977447, -44.918888075, 78.0650685987};
test_label[2755] = '{96.3573047515};
test_output[2755] = '{2.13293399321};
############ END DEBUG ############*/
test_input[22048:22055] = '{32'hc2a3297f, 32'hc28497c0, 32'h424dff7e, 32'h42026116, 32'hc20cafce, 32'hc2b65f4d, 32'hc25424cf, 32'h427d4630};
test_label[2756] = '{32'hc28497c0};
test_output[2756] = '{32'h43019d6c};
/*############ DEBUG ############
test_input[22048:22055] = '{-81.5810442169, -66.296387786, 51.4995057186, 32.5948108178, -35.1716826501, -91.1861378829, -53.035946823, 63.3185413242};
test_label[2756] = '{-66.296387786};
test_output[2756] = '{129.614936473};
############ END DEBUG ############*/
test_input[22056:22063] = '{32'h42a5af48, 32'h4225a186, 32'hc1b98c9f, 32'h42a4477b, 32'hc09da5f6, 32'h427b0765, 32'hc2175d0d, 32'hc243a180};
test_label[2757] = '{32'h4225a186};
test_output[2757] = '{32'h422758fa};
/*############ DEBUG ############
test_input[22056:22063] = '{82.8423489835, 41.4077366001, -23.1936635502, 82.1396088661, -4.92650910333, 62.7572226708, -37.840868842, -48.9077131547};
test_label[2757] = '{41.4077366001};
test_output[2757] = '{41.8368900611};
############ END DEBUG ############*/
test_input[22064:22071] = '{32'hc296b7d5, 32'hc286bd8e, 32'hc2c32687, 32'hc2c2248f, 32'h4259c927, 32'h42c5fb9e, 32'hc2bd5557, 32'h425fa0ea};
test_label[2758] = '{32'h4259c927};
test_output[2758] = '{32'h42322e15};
/*############ DEBUG ############
test_input[22064:22071] = '{-75.3590482967, -67.3702263293, -97.5752521687, -97.0713997833, 54.4464380334, 98.9914410449, -94.6666811915, 55.9071425157};
test_label[2758] = '{54.4464380334};
test_output[2758] = '{44.5450030115};
############ END DEBUG ############*/
test_input[22072:22079] = '{32'h42ad33e2, 32'h41bcc7ed, 32'hc2a3b2b9, 32'hbfcc1e09, 32'hc0ed1303, 32'h4205eb3f, 32'hc25c8876, 32'h429dd823};
test_label[2759] = '{32'hc25c8876};
test_output[2759] = '{32'h430dbc2d};
/*############ DEBUG ############
test_input[22072:22079] = '{86.6013301324, 23.5976194834, -81.8490643208, -1.59466654315, -7.40857074437, 33.4797326929, -55.1332637094, 78.9221442282};
test_label[2759] = '{-55.1332637094};
test_output[2759] = '{141.735056086};
############ END DEBUG ############*/
test_input[22080:22087] = '{32'h42c41616, 32'h426909c7, 32'hc267b51d, 32'h42b6372f, 32'h429fa1c7, 32'hc0a93b6e, 32'hc2bc21c2, 32'hc2b7dc35};
test_label[2760] = '{32'hc2b7dc35};
test_output[2760] = '{32'h433df966};
/*############ DEBUG ############
test_input[22080:22087] = '{98.0431400264, 58.2595498193, -57.9268674698, 91.1077780506, 79.8159704334, -5.28850445125, -94.0659322997, -91.9300936877};
test_label[2760] = '{-91.9300936877};
test_output[2760] = '{189.974206024};
############ END DEBUG ############*/
test_input[22088:22095] = '{32'hc2ba7792, 32'h42af5db5, 32'hc2716b59, 32'hc182dbff, 32'hc2a84e2c, 32'hc2943bfe, 32'h42783aa7, 32'h416e68f0};
test_label[2761] = '{32'h416e68f0};
test_output[2761] = '{32'h42919097};
/*############ DEBUG ############
test_input[22088:22095] = '{-93.2335374556, 87.6830215854, -60.3548318234, -16.3574201542, -84.1526810123, -74.117175179, 62.0572782236, 14.9006198404};
test_label[2761] = '{14.9006198404};
test_output[2761] = '{72.782401745};
############ END DEBUG ############*/
test_input[22096:22103] = '{32'hc1b684f4, 32'h42591585, 32'hc2485954, 32'hc181fca0, 32'hc2a37f2a, 32'h429b00ca, 32'h428eca21, 32'h42161d22};
test_label[2762] = '{32'h429b00ca};
test_output[2762] = '{32'h3b11d631};
/*############ DEBUG ############
test_input[22096:22103] = '{-22.8149194572, 54.2710161203, -50.0872361028, -16.2483513156, -81.7483670267, 77.5015389726, 71.3947842767, 37.5284507584};
test_label[2762] = '{77.5015389726};
test_output[2762] = '{0.00222529116521};
############ END DEBUG ############*/
test_input[22104:22111] = '{32'hc261a43d, 32'h4296937a, 32'hc2c0c8dd, 32'hc24c49d5, 32'h41baa908, 32'hc211ae13, 32'hc2722722, 32'hc09138a5};
test_label[2763] = '{32'h4296937a};
test_output[2763] = '{32'h80000000};
/*############ DEBUG ############
test_input[22104:22111] = '{-56.4103891499, 75.2880393153, -96.3923110024, -51.0721016334, 23.3325348374, -36.41999389, -60.5382146922, -4.53816479616};
test_label[2763] = '{75.2880393153};
test_output[2763] = '{-0.0};
############ END DEBUG ############*/
test_input[22112:22119] = '{32'hc1484a48, 32'hc20af620, 32'hc28f4d78, 32'hc0fb806e, 32'h4194d1fc, 32'h41f13933, 32'h42975d1b, 32'hc2b593ad};
test_label[2764] = '{32'h4194d1fc};
test_output[2764] = '{32'h42645137};
/*############ DEBUG ############
test_input[22112:22119] = '{-12.518134785, -34.7403570929, -71.6513059715, -7.85942721897, 18.6025322578, 30.1529298701, 75.6818449413, -90.788427908};
test_label[2764] = '{18.6025322578};
test_output[2764] = '{57.0793126834};
############ END DEBUG ############*/
test_input[22120:22127] = '{32'h42baa583, 32'h418a6590, 32'hc21e8000, 32'h41637dd5, 32'h428af3b1, 32'hc269c4da, 32'h42149f2a, 32'hc2867532};
test_label[2765] = '{32'h42baa583};
test_output[2765] = '{32'h2e416c20};
/*############ DEBUG ############
test_input[22120:22127] = '{93.3232637846, 17.2995913721, -39.6249982538, 14.2182211829, 69.4759584223, -58.4422394886, 37.155434729, -67.2288943261};
test_label[2765] = '{93.3232637846};
test_output[2765] = '{4.39791536531e-11};
############ END DEBUG ############*/
test_input[22128:22135] = '{32'hc26bc9ff, 32'hc1ef1504, 32'h41ade90d, 32'hc2a2c404, 32'h429df395, 32'h42902d9f, 32'h42c25476, 32'hbed98434};
test_label[2766] = '{32'h42c25476};
test_output[2766] = '{32'h3258c336};
/*############ DEBUG ############
test_input[22128:22135] = '{-58.9472625938, -29.8852618623, 21.7387951948, -81.3828401582, 78.9757423803, 72.0891072243, 97.1649648776, -0.424836766524};
test_label[2766] = '{97.1649648776};
test_output[2766] = '{1.26172403322e-08};
############ END DEBUG ############*/
test_input[22136:22143] = '{32'hbf3eb5e2, 32'h41a0de78, 32'hc29d34cd, 32'h416a6fb1, 32'h42bb3705, 32'hc2a983bc, 32'h419b42a4, 32'hc20213ff};
test_label[2767] = '{32'hbf3eb5e2};
test_output[2767] = '{32'h42bcb471};
/*############ DEBUG ############
test_input[22136:22143] = '{-0.744962811464, 20.1086268817, -78.6031302646, 14.652268352, 93.6074612803, -84.7572918627, 19.4075402481, -32.5195278627};
test_label[2767] = '{-0.744962811464};
test_output[2767] = '{94.3524240918};
############ END DEBUG ############*/
test_input[22144:22151] = '{32'h4240f3a0, 32'hc15dc087, 32'h424ff2c4, 32'h423247c3, 32'h424e180c, 32'h42a84b9f, 32'hc20831aa, 32'hc2b5011c};
test_label[2768] = '{32'hc2b5011c};
test_output[2768] = '{32'h432ea65d};
/*############ DEBUG ############
test_input[22144:22151] = '{48.2379155155, -13.8595036232, 51.9870754102, 44.5700803478, 51.5234849963, 84.1476953495, -34.0484997891, -90.5021634812};
test_label[2768] = '{-90.5021634812};
test_output[2768] = '{174.649858831};
############ END DEBUG ############*/
test_input[22152:22159] = '{32'hc049cbe6, 32'h42618f37, 32'hc295c31a, 32'h423b35bb, 32'h42449038, 32'h42c46d46, 32'hc2a6bdd3, 32'h422d3015};
test_label[2769] = '{32'h423b35bb};
test_output[2769] = '{32'h424da4d2};
/*############ DEBUG ############
test_input[22152:22159] = '{-3.15307004823, 56.3898586757, -74.8810562946, 46.8024693311, 49.1408392261, 98.2134282829, -83.3707490466, 43.2969564125};
test_label[2769] = '{46.8024693311};
test_output[2769] = '{51.4109589518};
############ END DEBUG ############*/
test_input[22160:22167] = '{32'h42318cfd, 32'h41b4adda, 32'hc27499af, 32'hc2ab3fa0, 32'h426c8373, 32'hc08bb1f9, 32'h4283612f, 32'h4046af6f};
test_label[2770] = '{32'h426c8373};
test_output[2770] = '{32'h40d202f3};
/*############ DEBUG ############
test_input[22160:22167] = '{44.3876829478, 22.5848888741, -61.1500829852, -85.6242695482, 59.1283675597, -4.36547539373, 65.6898147775, 3.10445765021};
test_label[2770] = '{59.1283675597};
test_output[2770] = '{6.56286005795};
############ END DEBUG ############*/
test_input[22168:22175] = '{32'hc21178c0, 32'hc1a93f98, 32'hc2940577, 32'h4260c2e2, 32'h42317145, 32'hc2c02b56, 32'h40a0f8f6, 32'hc2747a0e};
test_label[2771] = '{32'h4260c2e2};
test_output[2771] = '{32'h36f470e2};
/*############ DEBUG ############
test_input[22168:22175] = '{-36.3679197829, -21.1560511355, -74.0106742086, 56.1903153718, 44.3606132408, -96.084636828, 5.03039090925, -61.119193133};
test_label[2771] = '{56.1903153718};
test_output[2771] = '{7.28490780754e-06};
############ END DEBUG ############*/
test_input[22176:22183] = '{32'hc10209f1, 32'hc24c98fd, 32'h4257c383, 32'hc2b12134, 32'h41e023be, 32'hc2203486, 32'h406d4dac, 32'h40fea81b};
test_label[2772] = '{32'hc2203486};
test_output[2772] = '{32'h42bbfc05};
/*############ DEBUG ############
test_input[22176:22183] = '{-8.12742710385, -51.1494035352, 53.9409298551, -88.5648491736, 28.0174522178, -40.0512926283, 3.70786564027, 7.95802050706};
test_label[2772] = '{-40.0512926283};
test_output[2772] = '{93.9922224834};
############ END DEBUG ############*/
test_input[22184:22191] = '{32'hc1f8ec5f, 32'h42a1a9c3, 32'h4292c4a8, 32'hc22ac565, 32'hc28a9e84, 32'h428e8463, 32'hc2c2def1, 32'h41d1886b};
test_label[2773] = '{32'h4292c4a8};
test_output[2773] = '{32'h40ee5710};
/*############ DEBUG ############
test_input[22184:22191] = '{-31.1154153702, 80.8315694471, 73.3840941805, -42.6927662161, -69.3096025992, 71.2585662603, -97.4354355516, 26.1916108828};
test_label[2773] = '{73.3840941805};
test_output[2773] = '{7.44812754741};
############ END DEBUG ############*/
test_input[22192:22199] = '{32'hc182ecd4, 32'h42321e13, 32'h429dddc2, 32'hc2beb335, 32'hc270b645, 32'hc207651a, 32'hc1cd83ac, 32'h415be3e2};
test_label[2774] = '{32'hc2beb335};
test_output[2774] = '{32'h432e487c};
/*############ DEBUG ############
test_input[22192:22199] = '{-16.3656381843, 44.5293694512, 78.9331241641, -95.3500108957, -60.1779975281, -33.8487313848, -25.6892924354, 13.7431351317};
test_label[2774] = '{-95.3500108957};
test_output[2774] = '{174.28313506};
############ END DEBUG ############*/
test_input[22200:22207] = '{32'h406bed99, 32'h428c432f, 32'hc2b5408e, 32'hc20d80f5, 32'hc2191591, 32'h42762e31, 32'h42b32650, 32'hc27e1908};
test_label[2775] = '{32'h42762e31};
test_output[2775] = '{32'h41e03ce0};
/*############ DEBUG ############
test_input[22200:22207] = '{3.68637680202, 70.1312199068, -90.6260860356, -35.3759343787, -38.2710604407, 61.545107723, 89.5748316104, -63.5244439916};
test_label[2775] = '{61.545107723};
test_output[2775] = '{28.029723891};
############ END DEBUG ############*/
test_input[22208:22215] = '{32'h4279869a, 32'hbf7a0cc3, 32'h420a87ec, 32'hc1ff549d, 32'h41e2c278, 32'h42b5f266, 32'h4201b48e, 32'h4227b253};
test_label[2776] = '{32'h41e2c278};
test_output[2776] = '{32'h427a8391};
/*############ DEBUG ############
test_input[22208:22215] = '{62.3814468531, -0.976757223883, 34.6327352399, -31.9163156729, 28.3449559073, 90.9734378053, 32.4263235569, 41.9241437487};
test_label[2776] = '{28.3449559073};
test_output[2776] = '{62.628481898};
############ END DEBUG ############*/
test_input[22216:22223] = '{32'hc2bbdb34, 32'h423a0324, 32'h422d8352, 32'h4135607a, 32'hc297a968, 32'hc2862b9d, 32'h42c45881, 32'h42bed292};
test_label[2777] = '{32'h422d8352};
test_output[2777] = '{32'h425b6c6f};
/*############ DEBUG ############
test_input[22216:22223] = '{-93.9281286773, 46.5030689061, 43.3782416759, 11.3360541641, -75.8308688441, -67.0851838765, 98.1728576033, 95.411266716};
test_label[2777] = '{43.3782416759};
test_output[2777] = '{54.8558908397};
############ END DEBUG ############*/
test_input[22224:22231] = '{32'h42839a96, 32'h420a074a, 32'hc2c2da74, 32'hc2985ec3, 32'hc29dcf62, 32'hc2c1b05a, 32'hc12e68b9, 32'hc0fc7d40};
test_label[2778] = '{32'hc2c1b05a};
test_output[2778] = '{32'h4322a578};
/*############ DEBUG ############
test_input[22224:22231] = '{65.8019289362, 34.5071189816, -97.4266668951, -76.1850801245, -78.9050437595, -96.8444399894, -10.9005674872, -7.89028910482};
test_label[2778] = '{-96.8444399894};
test_output[2778] = '{162.646368926};
############ END DEBUG ############*/
test_input[22232:22239] = '{32'h42beefeb, 32'h425dc726, 32'h42bfc3b9, 32'hc26dfd7e, 32'h42339775, 32'hc26c2212, 32'h410bc396, 32'h4281d0a1};
test_label[2779] = '{32'h4281d0a1};
test_output[2779] = '{32'h41fbdbd3};
/*############ DEBUG ############
test_input[22232:22239] = '{95.4685864889, 55.444482014, 95.8822678911, -59.4975509306, 44.8979058158, -59.0332717589, 8.73525010779, 64.9074791834};
test_label[2779] = '{64.9074791834};
test_output[2779] = '{31.4823359102};
############ END DEBUG ############*/
test_input[22240:22247] = '{32'h42b54ca7, 32'h41aafa31, 32'h42993a9c, 32'hc2a62440, 32'hc243a513, 32'h4147b41f, 32'hc257ddc9, 32'hc1fe442c};
test_label[2780] = '{32'hc257ddc9};
test_output[2780] = '{32'h43109dc6};
/*############ DEBUG ############
test_input[22240:22247] = '{90.6497121555, 21.3721643257, 76.6144729337, -83.0707976789, -48.9112058272, 12.4814749981, -53.9665879128, -31.7832877823};
test_label[2780] = '{-53.9665879128};
test_output[2780] = '{144.616300871};
############ END DEBUG ############*/
test_input[22248:22255] = '{32'h40ab9bef, 32'hc17a7f2a, 32'h41b21da3, 32'hc235ac17, 32'h42100b87, 32'h41f11634, 32'hc26b3899, 32'h42990495};
test_label[2781] = '{32'h42100b87};
test_output[2781] = '{32'h4221fda3};
/*############ DEBUG ############
test_input[22248:22255] = '{5.36278478089, -15.6560454495, 22.2644717915, -45.4180574854, 36.0112567765, 30.1358407061, -58.8052711611, 76.5089504228};
test_label[2781] = '{36.0112567765};
test_output[2781] = '{40.4976936463};
############ END DEBUG ############*/
test_input[22256:22263] = '{32'h41935165, 32'hbf617434, 32'hc16a0fb4, 32'h41179679, 32'hc29de253, 32'hc25369b7, 32'hc27feb1f, 32'hc1b9964d};
test_label[2782] = '{32'hc16a0fb4};
test_output[2782] = '{32'h42042cc2};
/*############ DEBUG ############
test_input[22256:22263] = '{18.4147439181, -0.880679393758, -14.6288335058, 9.47423641937, -78.9420432312, -52.8532383755, -63.9796120627, -23.1983893951};
test_label[2782] = '{-14.6288335058};
test_output[2782] = '{33.0437083941};
############ END DEBUG ############*/
test_input[22264:22271] = '{32'h422013f8, 32'hc248fda0, 32'h42b49ba4, 32'hc0fcf7f5, 32'hc156f40a, 32'h414fd47d, 32'h420c1f15, 32'h4294fa81};
test_label[2783] = '{32'hc156f40a};
test_output[2783] = '{32'h42cf7a26};
/*############ DEBUG ############
test_input[22264:22271] = '{40.0195019745, -50.2476816989, 90.3039892093, -7.90526795428, -13.4345794839, 12.9893770833, 35.0303543686, 74.4892621497};
test_label[2783] = '{-13.4345794839};
test_output[2783] = '{103.738568829};
############ END DEBUG ############*/
test_input[22272:22279] = '{32'hc23b4b87, 32'h42a7555f, 32'h42865547, 32'h41f6aeed, 32'hc1f796f1, 32'hc18c59a6, 32'hc25294ec, 32'hc0f462c2};
test_label[2784] = '{32'hc0f462c2};
test_output[2784] = '{32'h42b69b8b};
/*############ DEBUG ############
test_input[22272:22279] = '{-46.8237562163, 83.6667423965, 67.1665562698, 30.8354139034, -30.9487026793, -17.5437744155, -52.6454305142, -7.63705546054};
test_label[2784] = '{-7.63705546054};
test_output[2784] = '{91.3037979253};
############ END DEBUG ############*/
test_input[22280:22287] = '{32'h4261f173, 32'hc0045bb3, 32'hc269bf00, 32'hc29dd3ba, 32'hc232a7e5, 32'hc1a25613, 32'h40d71a30, 32'hc264635f};
test_label[2785] = '{32'hc0045bb3};
test_output[2785] = '{32'h426a372f};
/*############ DEBUG ############
test_input[22280:22287] = '{56.4857914698, -2.06809687996, -58.4365218352, -78.9135285643, -44.6639586984, -20.2920282255, 6.72194675938, -57.0970423789};
test_label[2785] = '{-2.06809687996};
test_output[2785] = '{58.5538883497};
############ END DEBUG ############*/
test_input[22288:22295] = '{32'hc29f7f53, 32'hc2c2a142, 32'hc21326e5, 32'hc21e58e0, 32'h4191d035, 32'h42bd7989, 32'h42b2e6f1, 32'h4237c04c};
test_label[2786] = '{32'h4237c04c};
test_output[2786] = '{32'h424337f1};
/*############ DEBUG ############
test_input[22288:22295] = '{-79.7486822319, -97.3149595978, -36.7879841063, -39.5867930434, 18.226663394, 94.7373728401, 89.4510609184, 45.9377902324};
test_label[2786] = '{45.9377902324};
test_output[2786] = '{48.8046302359};
############ END DEBUG ############*/
test_input[22296:22303] = '{32'hc295523f, 32'h426fadc0, 32'hc2ae0189, 32'h41319619, 32'h42043073, 32'hc251d733, 32'h428adfb2, 32'hc26c0422};
test_label[2787] = '{32'h426fadc0};
test_output[2787] = '{32'h411846e0};
/*############ DEBUG ############
test_input[22296:22303] = '{-74.6606342907, 59.9196770311, -87.0029978958, 11.0991451014, 33.0473140223, -52.4601547996, 69.4369067712, -59.0040374933};
test_label[2787] = '{59.9196770311};
test_output[2787] = '{9.51730331054};
############ END DEBUG ############*/
test_input[22304:22311] = '{32'hc298b579, 32'h426277d7, 32'hc253be03, 32'hc2202dd8, 32'hc225c8cc, 32'h4288fbbf, 32'hc0566bb9, 32'h423a8b96};
test_label[2788] = '{32'hc298b579};
test_output[2788] = '{32'h4310d89c};
/*############ DEBUG ############
test_input[22304:22311] = '{-76.3544397083, 56.6170302402, -52.9355588227, -40.0447706525, -41.4460915512, 68.4916888441, -3.35032483675, 46.6363142269};
test_label[2788] = '{-76.3544397083};
test_output[2788] = '{144.846135517};
############ END DEBUG ############*/
test_input[22312:22319] = '{32'h424f0beb, 32'h42a2f704, 32'hc18e66ea, 32'h42365dc5, 32'hc241242c, 32'hc272f3dc, 32'hc26fcf59, 32'h4288489d};
test_label[2789] = '{32'h42a2f704};
test_output[2789] = '{32'h35d7ccb2};
/*############ DEBUG ############
test_input[22312:22319] = '{51.7616375351, 81.4824493336, -17.8002501583, 45.5915716017, -48.2853232435, -60.7381449938, -59.9524884367, 68.1418263188};
test_label[2789] = '{81.4824493336};
test_output[2789] = '{1.60783220686e-06};
############ END DEBUG ############*/
test_input[22320:22327] = '{32'hc202612a, 32'h405b2b90, 32'hc0f3ed18, 32'hc28d4a23, 32'h4297269c, 32'hc204bcce, 32'h4249124a, 32'h41f03106};
test_label[2790] = '{32'h4249124a};
test_output[2790] = '{32'h41ca75dc};
/*############ DEBUG ############
test_input[22320:22327] = '{-32.5948882804, 3.42453388605, -7.62269190552, -70.6448000022, 75.5754096334, -33.1843777723, 50.2678608668, 30.0239371625};
test_label[2790] = '{50.2678608668};
test_output[2790] = '{25.3075487666};
############ END DEBUG ############*/
test_input[22328:22335] = '{32'h42bea083, 32'h4244d503, 32'hc287addc, 32'hc2b1d701, 32'h424f9adb, 32'hc2ae1a88, 32'hc19f3421, 32'h42bbc880};
test_label[2791] = '{32'hc287addc};
test_output[2791] = '{32'h43235e84};
/*############ DEBUG ############
test_input[22328:22335] = '{95.3135032268, 49.2080181378, -67.8395678227, -88.9199300015, 51.9012277304, -87.0518179634, -19.9004544171, 93.8916047971};
test_label[2791] = '{-67.8395678227};
test_output[2791] = '{163.369194477};
############ END DEBUG ############*/
test_input[22336:22343] = '{32'hbfaf1bef, 32'h4049fe6e, 32'h42af6455, 32'hc1b344ff, 32'hc22704c9, 32'h423481f7, 32'hc254dfd5, 32'hc0cc06c2};
test_label[2792] = '{32'hc1b344ff};
test_output[2792] = '{32'h42dc3595};
/*############ DEBUG ############
test_input[22336:22343] = '{-1.36803997014, 3.15615413912, 87.6959626781, -22.4086893698, -41.7546723254, 45.1269172901, -53.2185857779, -6.37582488416};
test_label[2792] = '{-22.4086893698};
test_output[2792] = '{110.104652048};
############ END DEBUG ############*/
test_input[22344:22351] = '{32'hc13a6998, 32'h42597d7a, 32'h429f10ea, 32'hc2bb6726, 32'h407a3053, 32'hc1f3ddd6, 32'h421f96d1, 32'hc2a3a734};
test_label[2793] = '{32'hc1f3ddd6};
test_output[2793] = '{32'h42dc0860};
/*############ DEBUG ############
test_input[22344:22351] = '{-11.6507797899, 54.372536864, 79.5330352938, -93.7014619385, 3.90919938271, -30.4833187799, 39.8972811896, -81.8265654517};
test_label[2793] = '{-30.4833187799};
test_output[2793] = '{110.016354074};
############ END DEBUG ############*/
test_input[22352:22359] = '{32'h41e84a29, 32'hc1c3982b, 32'hc2a37ed7, 32'hc226fc58, 32'hc23cad69, 32'h4294598d, 32'hc2aad985, 32'hc283a0a3};
test_label[2794] = '{32'hc283a0a3};
test_output[2794] = '{32'h430bfd18};
/*############ DEBUG ############
test_input[22352:22359] = '{29.0362110867, -24.4493011474, -81.7477363605, -41.7464289436, -47.1693448806, 74.1749065, -85.4248394985, -65.8137419843};
test_label[2794] = '{-65.8137419843};
test_output[2794] = '{139.988648484};
############ END DEBUG ############*/
test_input[22360:22367] = '{32'h42a46f11, 32'h4068417a, 32'h406282a5, 32'h42839f4e, 32'hc0acb987, 32'hc1248a89, 32'h41e6ff7c, 32'h42bc548c};
test_label[2795] = '{32'hc0acb987};
test_output[2795] = '{32'h42c72025};
/*############ DEBUG ############
test_input[22360:22367] = '{82.2169254289, 3.62899643818, 3.53922398168, 65.811142366, -5.39764731483, -10.2838216705, 28.8747485381, 94.1651292845};
test_label[2795] = '{-5.39764731483};
test_output[2795] = '{99.5627830702};
############ END DEBUG ############*/
test_input[22368:22375] = '{32'hc2712bdd, 32'hc2c406bb, 32'hc278c4ab, 32'hc02cf75a, 32'hc2612d3a, 32'hc13ff1b4, 32'h3fd9d299, 32'h41362a53};
test_label[2796] = '{32'hc2c406bb};
test_output[2796] = '{32'h42dacc0e};
/*############ DEBUG ############
test_input[22368:22375] = '{-60.292837132, -98.0131450261, -62.19205725, -2.70259706211, -56.2941649723, -11.9965098553, 1.70173948099, 11.3853330924};
test_label[2796] = '{-98.0131450261};
test_output[2796] = '{109.398541175};
############ END DEBUG ############*/
test_input[22376:22383] = '{32'hc2b44055, 32'h426d483f, 32'hc2a5422c, 32'h427cac15, 32'hc1c70645, 32'hc2b1723f, 32'h42560b2c, 32'h427b7d11};
test_label[2797] = '{32'h426d483f};
test_output[2797] = '{32'h408d4e1f};
/*############ DEBUG ############
test_input[22376:22383] = '{-90.1256481384, 59.3205533005, -82.6292438987, 63.1680487887, -24.878061411, -88.7231393702, 53.5109092145, 62.8721332741};
test_label[2797] = '{59.3205533005};
test_output[2797] = '{4.41578630228};
############ END DEBUG ############*/
test_input[22384:22391] = '{32'hc1e57505, 32'hc1dd5e4f, 32'hc2228cd1, 32'h4284144b, 32'h40c7c8d0, 32'hc1a1e1ee, 32'h429bad2f, 32'h418f8f3a};
test_label[2798] = '{32'h429bad2f};
test_output[2798] = '{32'h36fc28d3};
/*############ DEBUG ############
test_input[22384:22391] = '{-28.6821390237, -27.6710482501, -40.6375155098, 66.0396358863, 6.24326335162, -20.2353171763, 77.8382499109, 17.9449347381};
test_label[2798] = '{77.8382499109};
test_output[2798] = '{7.51493802187e-06};
############ END DEBUG ############*/
test_input[22392:22399] = '{32'hc2af1f87, 32'hc221dffa, 32'hc29a0f68, 32'h4280c482, 32'h42a86df9, 32'hc2119e80, 32'hc261554d, 32'h4296fcea};
test_label[2799] = '{32'h42a86df9};
test_output[2799] = '{32'h392b1109};
/*############ DEBUG ############
test_input[22392:22399] = '{-87.5615769085, -40.4687285931, -77.0300932948, 64.3838073626, 84.2147941133, -36.4047853237, -56.333301816, 75.4939697089};
test_label[2799] = '{84.2147941133};
test_output[2799] = '{0.000163141764049};
############ END DEBUG ############*/
test_input[22400:22407] = '{32'hc1f44ecc, 32'h42278c86, 32'hc2843402, 32'h40cb7cd2, 32'hc28f03b6, 32'h422a41ea, 32'hc29f5cff, 32'h40c87230};
test_label[2800] = '{32'hc28f03b6};
test_output[2800] = '{32'h42e4f704};
/*############ DEBUG ############
test_input[22400:22407] = '{-30.538474273, 41.8872308185, -66.1015740126, 6.35898694581, -71.5072517024, 42.5643693551, -79.6816343565, 6.26393866889};
test_label[2800] = '{-71.5072517024};
test_output[2800] = '{114.482450906};
############ END DEBUG ############*/
test_input[22408:22415] = '{32'h41c94725, 32'h42513078, 32'h426c9577, 32'h40744e49, 32'h42771604, 32'h409646d2, 32'hc2a3eab0, 32'h410cb27f};
test_label[2801] = '{32'h410cb27f};
test_output[2801] = '{32'h4254310b};
/*############ DEBUG ############
test_input[22408:22415] = '{25.1597383027, 52.2973342855, 59.1459636066, 3.81727818045, 61.7715006023, 4.69614513187, -81.958371695, 8.79357810258};
test_label[2801] = '{8.79357810258};
test_output[2801] = '{53.0478940586};
############ END DEBUG ############*/
test_input[22416:22423] = '{32'h41dc9649, 32'h41d60969, 32'h42be19fb, 32'h41e00084, 32'hc2687cc0, 32'hc2914b70, 32'h4293752d, 32'h42b25af1};
test_label[2802] = '{32'h41dc9649};
test_output[2802] = '{32'h4286f5d9};
/*############ DEBUG ############
test_input[22416:22423] = '{27.573380711, 26.7545951365, 95.0507411574, 28.0002524854, -58.121825872, -72.6473406209, 73.7288617216, 89.1776163517};
test_label[2802] = '{27.573380711};
test_output[2802] = '{67.4801705611};
############ END DEBUG ############*/
test_input[22424:22431] = '{32'h42b8c290, 32'h42c070dc, 32'hc2357382, 32'h42a5e531, 32'h42396f30, 32'h4227f21b, 32'h41a3bcbd, 32'h427c01e2};
test_label[2803] = '{32'h427c01e2};
test_output[2803] = '{32'h4204f59a};
/*############ DEBUG ############
test_input[22424:22431] = '{92.3800029802, 96.2204270299, -45.362802081, 82.94764166, 46.3585806384, 41.9864325404, 20.4671576673, 63.0018391122};
test_label[2803] = '{63.0018391122};
test_output[2803] = '{33.2398465527};
############ END DEBUG ############*/
test_input[22432:22439] = '{32'h421aa94e, 32'hc113c207, 32'h42839105, 32'h4254e49d, 32'h42be231f, 32'h42ba0706, 32'hc26a5129, 32'h42abdcb0};
test_label[2804] = '{32'h42ba0706};
test_output[2804] = '{32'h400b3bac};
/*############ DEBUG ############
test_input[22432:22439] = '{38.6653384149, -9.23486948766, 65.7832420862, 53.2232562962, 95.0685987325, 93.013719107, -58.5792588495, 85.9310298047};
test_label[2804] = '{93.013719107};
test_output[2804] = '{2.17551707598};
############ END DEBUG ############*/
test_input[22440:22447] = '{32'hc1ad7fa7, 32'hc2bc9730, 32'hc266c684, 32'hc19721f6, 32'h3ecf5c5c, 32'hc1576a74, 32'h4208a40c, 32'hc2b10ae6};
test_label[2805] = '{32'hc1576a74};
test_output[2805] = '{32'h423e7ea9};
/*############ DEBUG ############
test_input[22440:22447] = '{-21.6873307301, -94.2952899871, -57.693862136, -18.8915827205, 0.405001508911, -13.4634899236, 34.1602007379, -88.5212861161};
test_label[2805] = '{-13.4634899236};
test_output[2805] = '{47.6236906615};
############ END DEBUG ############*/
test_input[22448:22455] = '{32'h4281dddc, 32'h424b66a5, 32'h42717068, 32'h4167f5c7, 32'hbf034cd5, 32'hc23ea143, 32'hbca8c6b3, 32'h4207b876};
test_label[2806] = '{32'h424b66a5};
test_output[2806] = '{32'h41617e58};
/*############ DEBUG ############
test_input[22448:22455] = '{64.9333153727, 50.8502388244, 60.3597719287, 14.4975044491, -0.512891111482, -47.657481149, -0.0206025593355, 33.9301391097};
test_label[2806] = '{50.8502388244};
test_output[2806] = '{14.0933457263};
############ END DEBUG ############*/
test_input[22456:22463] = '{32'hc0a584db, 32'hc26561ea, 32'hc27a7505, 32'hc0ced729, 32'hc16a5489, 32'hc2c7fa41, 32'hc1b271a4, 32'h421fd8ff};
test_label[2807] = '{32'hc16a5489};
test_output[2807] = '{32'h425a6e21};
/*############ DEBUG ############
test_input[22456:22463] = '{-5.17246792801, -57.3456201202, -62.614275761, -6.4637647439, -14.6456385244, -99.9887795953, -22.3054878833, 39.9619093996};
test_label[2807] = '{-14.6456385244};
test_output[2807] = '{54.6075479239};
############ END DEBUG ############*/
test_input[22464:22471] = '{32'hc2a96af7, 32'hc1d5ae0b, 32'h419d46b2, 32'h4206b74b, 32'h42ae5d69, 32'h41437708, 32'h4202a88f, 32'h42a696d3};
test_label[2808] = '{32'hc2a96af7};
test_output[2808] = '{32'h432be961};
/*############ DEBUG ############
test_input[22464:22471] = '{-84.708915646, -26.7099821572, 19.6595182829, 33.6789988906, 87.1824391383, 12.2165601772, 32.6646064992, 83.2945809063};
test_label[2808] = '{-84.708915646};
test_output[2808] = '{171.911636887};
############ END DEBUG ############*/
test_input[22472:22479] = '{32'h42a6bbe8, 32'h405fdf07, 32'h42a46696, 32'hc11a1029, 32'hc2b5ffb2, 32'h4296e8c3, 32'h4296717e, 32'hc226b3b5};
test_label[2809] = '{32'hc2b5ffb2};
test_output[2809] = '{32'h432ea355};
/*############ DEBUG ############
test_input[22472:22479] = '{83.3670067797, 3.49798755427, 82.200364598, -9.62894553363, -90.9994015417, 75.4546099121, 75.2216639588, -41.6754943841};
test_label[2809] = '{-90.9994015417};
test_output[2809] = '{174.63801216};
############ END DEBUG ############*/
test_input[22480:22487] = '{32'h4252468b, 32'h41a2bba3, 32'hc1203577, 32'h4038fb43, 32'h426505d4, 32'h3fa9c07c, 32'hc2789721, 32'h428b0662};
test_label[2810] = '{32'hc2789721};
test_output[2810] = '{32'h4303a8fa};
/*############ DEBUG ############
test_input[22480:22487] = '{52.568890458, 20.3416188915, -10.0130528928, 2.89033581853, 57.2556903763, 1.32618664162, -62.1475878022, 69.512467218};
test_label[2810] = '{-62.1475878022};
test_output[2810] = '{131.660059817};
############ END DEBUG ############*/
test_input[22488:22495] = '{32'h426d9451, 32'h4143c162, 32'hc157864c, 32'hc232bdaf, 32'hc119453b, 32'hc2bd5023, 32'h41d730fd, 32'hc13cf4af};
test_label[2811] = '{32'h41d730fd};
test_output[2811] = '{32'h4201fbd3};
/*############ DEBUG ############
test_input[22488:22495] = '{59.394841369, 12.2347128277, -13.4702875867, -44.6852364624, -9.57940170191, -94.6565184479, 26.8989197274, -11.8097368404};
test_label[2811] = '{26.8989197274};
test_output[2811] = '{32.4959216416};
############ END DEBUG ############*/
test_input[22496:22503] = '{32'hc2b60ea3, 32'h428309a8, 32'hc28203c2, 32'h41b06d0e, 32'h4149798d, 32'h42958001, 32'h42885991, 32'hc216760a};
test_label[2812] = '{32'hc216760a};
test_output[2812] = '{32'h42e0bbca};
/*############ DEBUG ############
test_input[22496:22503] = '{-91.028585274, 65.5188627688, -65.0073395152, 22.0532487185, 12.5921758554, 74.7500112018, 68.1749353592, -37.6152710843};
test_label[2812] = '{-37.6152710843};
test_output[2812] = '{112.366773814};
############ END DEBUG ############*/
test_input[22504:22511] = '{32'hc2823177, 32'hc28766c9, 32'hc293114e, 32'h4226fd4e, 32'h423dc4d5, 32'hc27dc23c, 32'h4269e9e0, 32'hc20c270a};
test_label[2813] = '{32'hc20c270a};
test_output[2813] = '{32'h42bb0877};
/*############ DEBUG ############
test_input[22504:22511] = '{-65.0966141354, -67.7007513793, -73.5337973272, 41.7473688501, 47.4422175061, -63.4396820044, 58.4783950923, -35.038124744};
test_label[2813] = '{-35.038124744};
test_output[2813] = '{93.5165359986};
############ END DEBUG ############*/
test_input[22512:22519] = '{32'h429c266a, 32'h427782a8, 32'hc2b03b28, 32'hc2835808, 32'h42140a05, 32'hc231824b, 32'hc267e319, 32'h422b4560};
test_label[2814] = '{32'h429c266a};
test_output[2814] = '{32'h33c65e76};
/*############ DEBUG ############
test_input[22512:22519] = '{78.0750271175, 61.8775934513, -88.1155359835, -65.6719385949, 37.0097834453, -44.3772392264, -57.9717762134, 42.8177493774};
test_label[2814] = '{78.0750271175};
test_output[2814] = '{9.23727599331e-08};
############ END DEBUG ############*/
test_input[22520:22527] = '{32'h4278e9f8, 32'h41a2db6a, 32'h40d3693e, 32'hc2bad71e, 32'hc2b914de, 32'h41af0df6, 32'h412581e8, 32'h428aea34};
test_label[2815] = '{32'hc2b914de};
test_output[2815] = '{32'h4321ffb9};
/*############ DEBUG ############
test_input[22520:22527] = '{62.2284867204, 20.357135743, 6.6065968545, -93.4201473892, -92.5407557082, 21.8818178044, 10.3442152858, 69.4574284627};
test_label[2815] = '{-92.5407557082};
test_output[2815] = '{161.998909196};
############ END DEBUG ############*/
test_input[22528:22535] = '{32'h40d97d19, 32'hc1cab47b, 32'hc269c6df, 32'h4218c120, 32'hc1c4214d, 32'h40d765f1, 32'hc2431a9f, 32'h414cb0a7};
test_label[2816] = '{32'hc1c4214d};
test_output[2816] = '{32'h427ad1c6};
/*############ DEBUG ############
test_input[22528:22535] = '{6.79652077388, -25.3381254361, -58.4442082993, 38.1885967793, -24.5162603223, 6.73119413122, -48.7759956616, 12.7931281512};
test_label[2816] = '{-24.5162603223};
test_output[2816] = '{62.7048571016};
############ END DEBUG ############*/
test_input[22536:22543] = '{32'hc283c651, 32'hbf31f0fd, 32'h40015ae7, 32'h42a34199, 32'hc2b7f5fa, 32'hc242b59b, 32'h42be2c52, 32'h4256e243};
test_label[2817] = '{32'hbf31f0fd};
test_output[2817] = '{32'h42bf9034};
/*############ DEBUG ############
test_input[22536:22543] = '{-65.8873381964, -0.695083458372, 2.02117329172, 81.6281211206, -91.9804209029, -48.677350688, 95.0865618182, 53.7209593113};
test_label[2817] = '{-0.695083458372};
test_output[2817] = '{95.7816467057};
############ END DEBUG ############*/
test_input[22544:22551] = '{32'h41eef9b4, 32'h429c67f2, 32'h42842576, 32'h41ba6946, 32'h407b940e, 32'hc225a468, 32'h41a2d70a, 32'hc26fc212};
test_label[2818] = '{32'h41eef9b4};
test_output[2818] = '{32'h4241530a};
/*############ DEBUG ############
test_input[22544:22551] = '{29.8719259258, 78.203015133, 66.0731624617, 23.3014031123, 3.93091157917, -41.4105514102, 20.3549997829, -59.9395201823};
test_label[2818] = '{29.8719259258};
test_output[2818] = '{48.3310946032};
############ END DEBUG ############*/
test_input[22552:22559] = '{32'h41f90e8d, 32'hc210f7d2, 32'hc222a5ad, 32'h428fbaf7, 32'hc1f302b5, 32'h4288c486, 32'h42be977b, 32'hc295919b};
test_label[2819] = '{32'h42be977b};
test_output[2819] = '{32'h2e9734d0};
/*############ DEBUG ############
test_input[22552:22559] = '{31.1321046572, -36.2420129978, -40.6617922446, 71.8651651885, -30.3763218056, 68.3838364905, 95.2958570804, -74.7843860371};
test_label[2819] = '{95.2958570804};
test_output[2819] = '{6.87606638318e-11};
############ END DEBUG ############*/
test_input[22560:22567] = '{32'hc26cd451, 32'h429b334e, 32'h425b6157, 32'h423aa93b, 32'hc2692e6e, 32'hc1fcfb0f, 32'hc190f241, 32'h42868112};
test_label[2820] = '{32'h429b334e};
test_output[2820] = '{32'h380670a2};
/*############ DEBUG ############
test_input[22560:22567] = '{-59.2073416664, 77.6002015671, 54.8450593493, 46.6652642769, -58.2953430849, -31.6225872724, -18.1182883084, 67.2520932755};
test_label[2820] = '{77.6002015671};
test_output[2820] = '{3.20529855099e-05};
############ END DEBUG ############*/
test_input[22568:22575] = '{32'h429ff6c5, 32'h41ce3e09, 32'h4226d01d, 32'hc0aeebd9, 32'hc2899bfb, 32'hc2b0f305, 32'hc1a1c406, 32'hc2862ba5};
test_label[2821] = '{32'hc0aeebd9};
test_output[2821] = '{32'h42aae582};
/*############ DEBUG ############
test_input[22568:22575] = '{79.9819680255, 25.7802906509, 41.7032347241, -5.4662899879, -68.8046456155, -88.474646911, -20.2207141229, -67.0852413357};
test_label[2821] = '{-5.4662899879};
test_output[2821] = '{85.4482580134};
############ END DEBUG ############*/
test_input[22576:22583] = '{32'hc28b0d9c, 32'hc2102613, 32'hc1b79ab2, 32'h417364ec, 32'h42c18832, 32'hc2835602, 32'h420d925d, 32'h428defe6};
test_label[2822] = '{32'h417364ec};
test_output[2822] = '{32'h42a31b94};
/*############ DEBUG ############
test_input[22576:22583] = '{-69.5265838259, -36.0371814568, -22.9505340062, 15.2121393422, 96.7660028329, -65.6679832899, 35.3929331617, 70.9685548565};
test_label[2822] = '{15.2121393422};
test_output[2822] = '{81.5538634908};
############ END DEBUG ############*/
test_input[22584:22591] = '{32'h3f51940a, 32'hc2824839, 32'hc21153cc, 32'hbf8962bc, 32'h426d6e35, 32'hc2089423, 32'hc1b9740f, 32'hc28b9e74};
test_label[2823] = '{32'hc21153cc};
test_output[2823] = '{32'h42bf6100};
/*############ DEBUG ############
test_input[22584:22591] = '{0.818665171296, -65.1410617023, -36.3318335947, -1.07332566783, 59.3576229561, -34.144666392, -23.1816687058, -69.8094774773};
test_label[2823] = '{-36.3318335947};
test_output[2823] = '{95.6894565508};
############ END DEBUG ############*/
test_input[22592:22599] = '{32'hc17cf815, 32'h4289fb70, 32'hc0c3d6aa, 32'hc0a1f07f, 32'hc134d54b, 32'hc16e4904, 32'hc20985cf, 32'h41f78f13};
test_label[2824] = '{32'hc17cf815};
test_output[2824] = '{32'h42a99a73};
/*############ DEBUG ############
test_input[22592:22599] = '{-15.8105664343, 68.9910884397, -6.11995422496, -5.06060728508, -11.3020738656, -14.8928261499, -34.3806733497, 30.9448610949};
test_label[2824] = '{-15.8105664343};
test_output[2824] = '{84.801654874};
############ END DEBUG ############*/
test_input[22600:22607] = '{32'h42012ce2, 32'hc26eef99, 32'hc28fe027, 32'h420fe886, 32'h4095f28a, 32'h42644352, 32'h42c12fbc, 32'h428ef035};
test_label[2825] = '{32'h420fe886};
test_output[2825] = '{32'h427276f3};
/*############ DEBUG ############
test_input[22600:22607] = '{32.293830496, -59.733981984, -71.93779898, 35.9770719566, 4.68585678012, 57.0657406551, 96.5932343581, 71.4691534273};
test_label[2825] = '{35.9770719566};
test_output[2825] = '{60.6161624015};
############ END DEBUG ############*/
test_input[22608:22615] = '{32'hc206a750, 32'hc27852b1, 32'h42af265b, 32'hc2babd1e, 32'hc2084714, 32'hc274abfd, 32'h41283acf, 32'hc2c01ccb};
test_label[2826] = '{32'hc27852b1};
test_output[2826] = '{32'h4315a7da};
/*############ DEBUG ############
test_input[22608:22615] = '{-33.6633915741, -62.0807550711, 87.5749160681, -93.3693705733, -34.0694112716, -61.1679568968, 10.5143578795, -96.0562332961};
test_label[2826] = '{-62.0807550711};
test_output[2826] = '{149.655671139};
############ END DEBUG ############*/
test_input[22616:22623] = '{32'h42482630, 32'h425349cd, 32'h42936f0c, 32'h42235483, 32'hc1098855, 32'h422bf501, 32'h408f0f54, 32'h41d97c61};
test_label[2827] = '{32'hc1098855};
test_output[2827] = '{32'h42a4a017};
/*############ DEBUG ############
test_input[22616:22623] = '{50.0372919115, 52.8220726085, 73.7168918265, 40.8325300703, -8.59578433441, 42.9892633075, 4.47062132587, 27.1857311752};
test_label[2827] = '{-8.59578433441};
test_output[2827] = '{82.3126761618};
############ END DEBUG ############*/
test_input[22624:22631] = '{32'hc286a86e, 32'h4282c2b6, 32'h42a60389, 32'hc2154816, 32'h41eb9cac, 32'hc25d403b, 32'hc20832cd, 32'hc07e997d};
test_label[2828] = '{32'hc2154816};
test_output[2828] = '{32'h42f0a794};
/*############ DEBUG ############
test_input[22624:22631] = '{-67.3289605592, 65.3802913591, 83.0069032962, -37.320395931, 29.4515005302, -55.312724279, -34.0496087139, -3.97811811593};
test_label[2828] = '{-37.320395931};
test_output[2828] = '{120.327299249};
############ END DEBUG ############*/
test_input[22632:22639] = '{32'h425d51a3, 32'h4005bbce, 32'h42b110c6, 32'h41b9e3b3, 32'hc2491e63, 32'h3fc8eb2d, 32'hc2be77f3, 32'h42675459};
test_label[2829] = '{32'h4005bbce};
test_output[2829] = '{32'h42ace2e8};
/*############ DEBUG ############
test_input[22632:22639] = '{55.3297229771, 2.08958780514, 88.5327625675, 23.2361815257, -50.2796737648, 1.56967696336, -95.2342782669, 57.8323710856};
test_label[2829] = '{2.08958780514};
test_output[2829] = '{86.4431747624};
############ END DEBUG ############*/
test_input[22640:22647] = '{32'hbf2f2687, 32'h4025a360, 32'h4137f49a, 32'hc12b583a, 32'h4294d6f3, 32'h4263c37c, 32'h4236c47c, 32'h42a7aa98};
test_label[2830] = '{32'h4263c37c};
test_output[2830] = '{32'h41d72390};
/*############ DEBUG ############
test_input[22640:22647] = '{-0.684181649595, 2.58809665619, 11.4972167335, -10.7090395977, 74.4198246291, 56.9409044384, 45.6918785702, 83.8331871386};
test_label[2830] = '{56.9409044384};
test_output[2830] = '{26.8923643229};
############ END DEBUG ############*/
test_input[22648:22655] = '{32'hc2a3724c, 32'hc293f118, 32'hc221dc64, 32'h42510e66, 32'hc2a6a1f1, 32'h417104ba, 32'hc2baa366, 32'hc0da655d};
test_label[2831] = '{32'hc0da655d};
test_output[2831] = '{32'h426c5b12};
/*############ DEBUG ############
test_input[22648:22655] = '{-81.7232397112, -73.9708870409, -40.4652238778, 52.2640606716, -83.3162953742, 15.0636541319, -93.3191396329, -6.82487344399};
test_label[2831] = '{-6.82487344399};
test_output[2831] = '{59.0889341155};
############ END DEBUG ############*/
test_input[22656:22663] = '{32'h41b6e7f0, 32'h420d2604, 32'h4129542e, 32'hc21501b0, 32'hc2adfc17, 32'hc19f2109, 32'hc1cb3997, 32'hc2817cb4};
test_label[2832] = '{32'hc2817cb4};
test_output[2832] = '{32'h42c80fb7};
/*############ DEBUG ############
test_input[22656:22663] = '{22.8632506492, 35.2871250858, 10.5830518756, -37.2516491443, -86.9923637115, -19.8911304621, -25.403120702, -64.7435621519};
test_label[2832] = '{-64.7435621519};
test_output[2832] = '{100.030691259};
############ END DEBUG ############*/
test_input[22664:22671] = '{32'hc1ab045e, 32'hc261bf39, 32'h413874fc, 32'h42811e8d, 32'h42661af5, 32'h424af3ce, 32'h40225c3d, 32'hc27f0b56};
test_label[2833] = '{32'h424af3ce};
test_output[2833] = '{32'h415d28ce};
/*############ DEBUG ############
test_input[22664:22671] = '{-21.3771316096, -56.4367406602, 11.5285609166, 64.5596698146, 57.5263254168, 50.7380905838, 2.53687982109, -63.7610708691};
test_label[2833] = '{50.7380905838};
test_output[2833] = '{13.8224618124};
############ END DEBUG ############*/
test_input[22672:22679] = '{32'hc23e2528, 32'hc084dd21, 32'h42237f12, 32'h42118bfb, 32'hc2113948, 32'h41111151, 32'h3fa60f0c, 32'h41ee77ef};
test_label[2834] = '{32'h3fa60f0c};
test_output[2834] = '{32'h421e5a12};
/*############ DEBUG ############
test_input[22672:22679] = '{-47.5362851152, -4.15199331229, 40.8740916648, 36.3866988878, -36.3059385896, 9.0667279911, 1.29733419095, 29.8085611166};
test_label[2834] = '{1.29733419095};
test_output[2834] = '{39.5879600688};
############ END DEBUG ############*/
test_input[22680:22687] = '{32'h41920219, 32'hc1b6118f, 32'hc289c1a3, 32'hc22609da, 32'h42c446ff, 32'h42a6e530, 32'h41af8905, 32'hc2028e39};
test_label[2835] = '{32'h41920219};
test_output[2835] = '{32'h429fc679};
/*############ DEBUG ############
test_input[22680:22687] = '{18.2510238271, -22.7585731863, -68.8781989467, -41.5096195508, 98.1386637371, 83.4476287528, 21.9419042794, -32.6388911223};
test_label[2835] = '{18.2510238271};
test_output[2835] = '{79.8876403266};
############ END DEBUG ############*/
test_input[22688:22695] = '{32'h40dac976, 32'hc2b90396, 32'h412957b3, 32'h424caf03, 32'hc29f121d, 32'h42b48b39, 32'h42535a6d, 32'hc116c242};
test_label[2836] = '{32'h412957b3};
test_output[2836] = '{32'h429f6043};
/*############ DEBUG ############
test_input[22688:22695] = '{6.83709253862, -92.5070018603, 10.5839105948, 51.1709116925, -79.535375915, 90.2719209097, 52.8383059345, -9.42242596233};
test_label[2836] = '{10.5839105948};
test_output[2836] = '{79.6880103149};
############ END DEBUG ############*/
test_input[22696:22703] = '{32'hc221c589, 32'hc2336c2c, 32'h41c06f22, 32'hc2a59cd0, 32'h42c25789, 32'hc28a7382, 32'hc0e31616, 32'h42c42a43};
test_label[2837] = '{32'h42c25789};
test_output[2837] = '{32'h3f9fec44};
/*############ DEBUG ############
test_input[22696:22703] = '{-40.4429056918, -44.8556382949, 24.0542643689, -82.8062750469, 97.1709651846, -69.2256010226, -7.09644597736, 98.082541413};
test_label[2837] = '{97.1709651846};
test_output[2837] = '{1.24939773556};
############ END DEBUG ############*/
test_input[22704:22711] = '{32'hc22980ea, 32'hc10ef8d6, 32'h42251d7d, 32'h42aabb9f, 32'h4112c8f9, 32'hc21bb71f, 32'h4221f6a4, 32'hc2848160};
test_label[2838] = '{32'h42251d7d};
test_output[2838] = '{32'h423059c2};
/*############ DEBUG ############
test_input[22704:22711] = '{-42.3758938217, -8.93575118962, 41.2787958928, 85.3664489648, 9.17406558075, -38.9288297542, 40.4908610099, -66.252687862};
test_label[2838] = '{41.2787958928};
test_output[2838] = '{44.087653072};
############ END DEBUG ############*/
test_input[22712:22719] = '{32'hc2b0f8de, 32'hc24efadd, 32'hc23ef320, 32'hc2099abc, 32'hc268f136, 32'hc131697e, 32'hc1c7125a, 32'hc23593de};
test_label[2839] = '{32'hc2b0f8de};
test_output[2839] = '{32'h429acbae};
/*############ DEBUG ############
test_input[22712:22719] = '{-88.4860665943, -51.7449844725, -47.7374262925, -34.401109451, -58.2355588917, -11.0882548437, -24.8839616159, -45.3944004271};
test_label[2839] = '{-88.4860665943};
test_output[2839] = '{77.3978127707};
############ END DEBUG ############*/
test_input[22720:22727] = '{32'hc21040fc, 32'h41be168b, 32'h428197ae, 32'h41ff8b06, 32'h42a311b1, 32'h427e0c99, 32'h41ec3169, 32'hc19de053};
test_label[2840] = '{32'h428197ae};
test_output[2840] = '{32'h4185e80b};
/*############ DEBUG ############
test_input[22720:22727] = '{-36.0634607825, 23.7610080397, 64.7962488285, 31.9428824319, 81.5345502823, 63.5123040366, 29.5241254519, -19.7345326555};
test_label[2840] = '{64.7962488285};
test_output[2840] = '{16.7383015224};
############ END DEBUG ############*/
test_input[22728:22735] = '{32'h4220da85, 32'h418332ea, 32'h4177bd2f, 32'h429111b2, 32'hc288da43, 32'hc23b5448, 32'hc260d8dc, 32'hc27e6f85};
test_label[2841] = '{32'h429111b2};
test_output[2841] = '{32'h28260000};
/*############ DEBUG ############
test_input[22728:22735] = '{40.2133967787, 16.3998598776, 15.4836872243, 72.5345621102, -68.4262919964, -46.8323070098, -56.2117762951, -63.6089066012};
test_label[2841] = '{72.5345621102};
test_output[2841] = '{9.21485110439e-15};
############ END DEBUG ############*/
test_input[22736:22743] = '{32'hc28930fa, 32'h41cb795b, 32'h427978fc, 32'hc285e977, 32'h42aa1d2c, 32'h42921dd6, 32'hc22b00b5, 32'hc1e18840};
test_label[2842] = '{32'h427978fc};
test_output[2842] = '{32'h41b582bb};
/*############ DEBUG ############
test_input[22736:22743] = '{-68.59565389, 25.4342558443, 62.3681484626, -66.9559871154, 85.0569754386, 73.0582766234, -42.7506896867, -28.1915287071};
test_label[2842] = '{62.3681484626};
test_output[2842] = '{22.6888331283};
############ END DEBUG ############*/
test_input[22744:22751] = '{32'h4287b36c, 32'hc0e30880, 32'h427283fd, 32'h4284c254, 32'h414c7453, 32'hc2bdcef1, 32'h422c5e5a, 32'hbfbc6d78};
test_label[2843] = '{32'h427283fd};
test_output[2843] = '{32'h40edb9bf};
/*############ DEBUG ############
test_input[22744:22751] = '{67.8504354725, -7.09478778697, 60.6288932284, 66.3795493689, 12.7783994795, -94.9041812273, 43.0921383927, -1.47209075562};
test_label[2843] = '{60.6288932284};
test_output[2843] = '{7.42892424206};
############ END DEBUG ############*/
test_input[22752:22759] = '{32'hc2c4ab09, 32'h428851a4, 32'hc1b82e35, 32'h42b9fa74, 32'hc294e86d, 32'h40c3dc85, 32'h423eb645, 32'hc2aa5f99};
test_label[2844] = '{32'h428851a4};
test_output[2844] = '{32'h41c6a33d};
/*############ DEBUG ############
test_input[22752:22759] = '{-98.3340498904, 68.1594578651, -23.0225626934, 92.9891638146, -74.4539573248, 6.12066906932, 47.6779970434, -85.186717786};
test_label[2844] = '{68.1594578651};
test_output[2844] = '{24.8297059496};
############ END DEBUG ############*/
test_input[22760:22767] = '{32'hc1908438, 32'h42c33007, 32'hc1fba862, 32'hc1bee8ff, 32'h41e7814f, 32'h41ae585d, 32'hc200fcc5, 32'hc19be3db};
test_label[2845] = '{32'h41ae585d};
test_output[2845] = '{32'h429799f0};
/*############ DEBUG ############
test_input[22760:22767] = '{-18.0645606977, 97.5938029287, -31.4572176085, -23.8637667947, 28.9381383416, 21.793147042, -32.2468466542, -19.4862569505};
test_label[2845] = '{21.793147042};
test_output[2845] = '{75.8006558868};
############ END DEBUG ############*/
test_input[22768:22775] = '{32'hc2b923fb, 32'hc1906070, 32'h419ff18b, 32'hc2a91540, 32'hc17f8747, 32'hc1fa2015, 32'hc1328a64, 32'h42c7cea6};
test_label[2846] = '{32'hc1328a64};
test_output[2846] = '{32'h42de1ff3};
/*############ DEBUG ############
test_input[22768:22775] = '{-92.5702752101, -18.0470879059, 19.9929412037, -84.5415064994, -15.970526862, -31.2656651693, -11.1587871027, 99.9036118678};
test_label[2846] = '{-11.1587871027};
test_output[2846] = '{111.06239897};
############ END DEBUG ############*/
test_input[22776:22783] = '{32'h40849192, 32'h4290a5d8, 32'h42579c59, 32'hc29e03ca, 32'hc2848759, 32'h425df7d3, 32'hc1bcc279, 32'h42bd9f49};
test_label[2847] = '{32'h4290a5d8};
test_output[2847] = '{32'h41b3e5c4};
/*############ DEBUG ############
test_input[22776:22783] = '{4.14276960921, 72.3239156443, 53.902684077, -79.0073998637, -66.2643515827, 55.4920165759, -23.5949571406, 94.8111051161};
test_label[2847] = '{72.3239156443};
test_output[2847] = '{22.487189472};
############ END DEBUG ############*/
test_input[22784:22791] = '{32'hc25fcc8b, 32'hc288d7a9, 32'hc22439d1, 32'hc1befa99, 32'h42a46640, 32'hc1acdcd1, 32'hc298f60b, 32'h42164a77};
test_label[2848] = '{32'hc298f60b};
test_output[2848] = '{32'h431eae26};
/*############ DEBUG ############
test_input[22784:22791] = '{-55.949747687, -68.4212141618, -41.0564605211, -23.8723615993, 82.1997107512, -21.6078204759, -76.4805561688, 37.5727210632};
test_label[2848] = '{-76.4805561688};
test_output[2848] = '{158.68026692};
############ END DEBUG ############*/
test_input[22792:22799] = '{32'h429a73b5, 32'h42b44f0c, 32'hc25bbea8, 32'hc03bafb6, 32'h4253ed88, 32'hc25d9bd5, 32'hc292a664, 32'hc24622e5};
test_label[2849] = '{32'hc24622e5};
test_output[2849] = '{32'h430bb040};
/*############ DEBUG ############
test_input[22792:22799] = '{77.2259910574, 90.1543899748, -54.9361879696, -2.93259947359, 52.9819625082, -55.4021804145, -73.324983204, -49.5340769307};
test_label[2849] = '{-49.5340769307};
test_output[2849] = '{139.688469334};
############ END DEBUG ############*/
test_input[22800:22807] = '{32'h4245620a, 32'h426c38d9, 32'hc21bfcc0, 32'hc2c1e12d, 32'hc1d10421, 32'hc288cfb4, 32'hc1984eb1, 32'hc2246e25};
test_label[2850] = '{32'hc1984eb1};
test_output[2850] = '{32'h429c3021};
/*############ DEBUG ############
test_input[22800:22807] = '{49.3457402242, 59.0555155985, -38.9968265888, -96.9398000322, -26.1270169827, -68.4056695494, -19.0384228349, -41.107562448};
test_label[2850] = '{-19.0384228349};
test_output[2850] = '{78.0939991189};
############ END DEBUG ############*/
test_input[22808:22815] = '{32'h42c0e9e0, 32'hc1699afa, 32'hc2362956, 32'h41d259fe, 32'hc299a903, 32'h426e6e8e, 32'hc28c44e8, 32'h41ea2094};
test_label[2851] = '{32'h41d259fe};
test_output[2851] = '{32'h428c5361};
/*############ DEBUG ############
test_input[22808:22815] = '{96.45678995, -14.6003356969, -45.5403665501, 26.2939412036, -76.830100151, 59.6079631462, -70.1345816739, 29.2659069763};
test_label[2851] = '{26.2939412036};
test_output[2851] = '{70.1628487463};
############ END DEBUG ############*/
test_input[22816:22823] = '{32'h40820203, 32'hc231f3b1, 32'h4295c86f, 32'h41c4569b, 32'h411feca5, 32'hbf8a8a35, 32'hc28f9ad9, 32'hc2847c42};
test_label[2852] = '{32'hc2847c42};
test_output[2852] = '{32'h430d2259};
/*############ DEBUG ############
test_input[22816:22823] = '{4.06274571918, -44.4879807127, 74.8914738595, 24.5422885971, 9.99527456128, -1.08234272083, -71.8024352261, -66.2426907768};
test_label[2852] = '{-66.2426907768};
test_output[2852] = '{141.134164636};
############ END DEBUG ############*/
test_input[22824:22831] = '{32'h4293243d, 32'h41afed6e, 32'h41aa096f, 32'h428a9aad, 32'h428a6b5b, 32'hc247dcb6, 32'hc2805914, 32'hc0ccbbbc};
test_label[2853] = '{32'h428a6b5b};
test_output[2853] = '{32'h408c6688};
/*############ DEBUG ############
test_input[22824:22831] = '{73.5707780765, 21.9909324886, 21.2546066263, 69.3021046182, 69.2096749942, -49.965539356, -64.1739838405, -6.39791666674};
test_label[2853] = '{69.2096749942};
test_output[2853] = '{4.38751581721};
############ END DEBUG ############*/
test_input[22832:22839] = '{32'hc27d2e4b, 32'hc0bd987b, 32'hc29a8ddb, 32'hc11db526, 32'hc274dd21, 32'hc2af7558, 32'h42b96288, 32'h40ffd340};
test_label[2854] = '{32'hc274dd21};
test_output[2854] = '{32'h4319e88c};
/*############ DEBUG ############
test_input[22832:22839] = '{-63.2952090374, -5.92486335057, -77.2770609485, -9.85672526427, -61.2159469789, -87.7291877524, 92.6924430535, 7.9945374209};
test_label[2854] = '{-61.2159469789};
test_output[2854] = '{153.908390032};
############ END DEBUG ############*/
test_input[22840:22847] = '{32'h40e075e6, 32'hc260cd61, 32'hc2929a2c, 32'hc244340e, 32'h429d462a, 32'h41ad2423, 32'hc28b9b32, 32'h423e21ff};
test_label[2855] = '{32'hc260cd61};
test_output[2855] = '{32'h4306d66d};
/*############ DEBUG ############
test_input[22840:22847] = '{7.01439194863, -56.2005653866, -73.3011141719, -49.0508330841, 78.6370421692, 21.6426455232, -69.80311529, 47.533200643};
test_label[2855] = '{-56.2005653866};
test_output[2855] = '{134.837607556};
############ END DEBUG ############*/
test_input[22848:22855] = '{32'hc29eb9d1, 32'hc200dd69, 32'hc11738e8, 32'h42601291, 32'h41b633eb, 32'hc19b6c99, 32'hc2b66b17, 32'hc1bb9521};
test_label[2856] = '{32'hc2b66b17};
test_output[2856] = '{32'h43133a30};
/*############ DEBUG ############
test_input[22848:22855] = '{-79.3629194697, -32.2162189902, -9.4513935853, 56.0181327356, 22.7753508909, -19.4280264556, -91.2091565971, -23.4478163551};
test_label[2856] = '{-91.2091565971};
test_output[2856] = '{147.227289333};
############ END DEBUG ############*/
test_input[22856:22863] = '{32'h421b4acc, 32'hc0801c5f, 32'hc2af9448, 32'h3eda6b6b, 32'hc248c406, 32'hc0f467ef, 32'h4233caf0, 32'hc24e5678};
test_label[2857] = '{32'hc0801c5f};
test_output[2857] = '{32'h4243d0b9};
/*############ DEBUG ############
test_input[22856:22863] = '{38.8230429537, -4.00346321883, -87.7896110882, 0.426600785186, -50.1914277631, -7.63768731116, 44.9481825781, -51.5844428182};
test_label[2857] = '{-4.00346321883};
test_output[2857] = '{48.9538305943};
############ END DEBUG ############*/
test_input[22864:22871] = '{32'hc2a4116c, 32'h422eb21f, 32'hc27e20be, 32'h41e73690, 32'h42486c0d, 32'h40d7bf41, 32'h42815dee, 32'hc280efc7};
test_label[2858] = '{32'h422eb21f};
test_output[2858] = '{32'h41a8137a};
/*############ DEBUG ############
test_input[22864:22871] = '{-82.0340288768, 43.6739456661, -63.5319755429, 28.9016427319, 50.1055176726, 6.74209647973, 64.683456087, -64.4683189159};
test_label[2858] = '{43.6739456661};
test_output[2858] = '{21.0095108881};
############ END DEBUG ############*/
test_input[22872:22879] = '{32'h3fa5afd8, 32'hc269c98d, 32'hc295b31d, 32'hc1b48981, 32'hc2abf837, 32'hc28c31a9, 32'hc242f596, 32'hc1c88d8b};
test_label[2859] = '{32'hc1c88d8b};
test_output[2859] = '{32'h41d2e889};
/*############ DEBUG ############
test_input[22872:22879] = '{1.29442885578, -58.4468257388, -74.8498325566, -22.5671401965, -85.9847916197, -70.0969931178, -48.7398313247, -25.069113652};
test_label[2859] = '{-25.069113652};
test_output[2859] = '{26.3635425079};
############ END DEBUG ############*/
test_input[22880:22887] = '{32'h41246e76, 32'hc2348d00, 32'hc0026f02, 32'h421894a1, 32'h3fd864f8, 32'h429c7f0e, 32'h428da168, 32'hc11e8e1f};
test_label[2860] = '{32'hc0026f02};
test_output[2860] = '{32'h42a092d3};
/*############ DEBUG ############
test_input[22880:22887] = '{10.276968179, -45.1376948661, -2.03802526267, 38.1451465442, 1.69058132906, 78.2481509636, 70.8152456794, -9.90969791279};
test_label[2860] = '{-2.03802526267};
test_output[2860] = '{80.286767518};
############ END DEBUG ############*/
test_input[22888:22895] = '{32'h4255ad1e, 32'h415c025e, 32'hc1fb81f6, 32'hc20c124c, 32'hc20237f0, 32'hc107eb2b, 32'hc191d384, 32'h42c681bf};
test_label[2861] = '{32'h4255ad1e};
test_output[2861] = '{32'h42375660};
/*############ DEBUG ############
test_input[22888:22895] = '{53.4190584914, 13.7505776263, -31.4384582042, -35.0178676597, -32.5546269565, -8.49491452412, -18.2282782253, 99.2534076821};
test_label[2861] = '{53.4190584914};
test_output[2861] = '{45.8343491907};
############ END DEBUG ############*/
test_input[22896:22903] = '{32'h41d1f7da, 32'h42c21299, 32'h42928eaf, 32'h4243ba37, 32'hc23009a9, 32'h42b0e07c, 32'h422131f4, 32'hc2c1a99f};
test_label[2862] = '{32'h4243ba37};
test_output[2862] = '{32'h42406b2b};
/*############ DEBUG ############
test_input[22896:22903] = '{26.2460205059, 97.0363244389, 73.2786779087, 48.9318513998, -44.0094347817, 88.4384471857, 40.2987839064, -96.8312901624};
test_label[2862] = '{48.9318513998};
test_output[2862] = '{48.1046575191};
############ END DEBUG ############*/
test_input[22904:22911] = '{32'h42c5be56, 32'hc236893e, 32'h41c2965f, 32'hc2ab0b0a, 32'h4211acf7, 32'hc21383be, 32'hc0eb892a, 32'h42422527};
test_label[2863] = '{32'h42422527};
test_output[2863] = '{32'h42495785};
/*############ DEBUG ############
test_input[22904:22911] = '{98.8717517583, -45.6340266562, 24.3234237384, -85.5215634672, 36.4189094918, -36.8786532635, -7.36049374385, 48.5362822866};
test_label[2863] = '{48.5362822866};
test_output[2863] = '{50.3354694717};
############ END DEBUG ############*/
test_input[22912:22919] = '{32'h42be93b5, 32'hc23fa11d, 32'h4158db68, 32'hc28ace0d, 32'hc223b228, 32'hc2bc3769, 32'h42846ab8, 32'hc2b22643};
test_label[2864] = '{32'hc2bc3769};
test_output[2864] = '{32'h433d658f};
/*############ DEBUG ############
test_input[22912:22919] = '{95.2884885611, -47.9073355398, 13.5535658246, -69.4024422995, -40.9239795106, -94.1082221206, 66.2084354485, -89.0747316504};
test_label[2864] = '{-94.1082221206};
test_output[2864] = '{189.396710682};
############ END DEBUG ############*/
test_input[22920:22927] = '{32'hc289864e, 32'h427f6d29, 32'h41ce439c, 32'hc28cfd65, 32'h413231fb, 32'hc279a3e5, 32'hbe834719, 32'h41693eba};
test_label[2865] = '{32'hc279a3e5};
test_output[2865] = '{32'h42fc8887};
/*############ DEBUG ############
test_input[22920:22927] = '{-68.7623144688, 63.8566029404, 25.7830115131, -70.4949107532, 11.1372025164, -62.4100539241, -0.256401807509, 14.5778144919};
test_label[2865] = '{-62.4100539241};
test_output[2865] = '{126.266656865};
############ END DEBUG ############*/
test_input[22928:22935] = '{32'h42b8ab20, 32'h40591ddc, 32'hc2162865, 32'hc1572713, 32'hc2470dde, 32'h4227bb06, 32'hc28ce9b5, 32'hbfebd208};
test_label[2866] = '{32'hc28ce9b5};
test_output[2866] = '{32'h4322ca6b};
/*############ DEBUG ############
test_input[22928:22935] = '{92.3342288129, 3.3924473694, -37.5394483307, -13.4470398786, -49.7635407245, 41.932639915, -70.4564590517, -1.84234717822};
test_label[2866] = '{-70.4564590517};
test_output[2866] = '{162.790687865};
############ END DEBUG ############*/
test_input[22936:22943] = '{32'hc295076d, 32'h422d3c32, 32'hc25113b7, 32'h4258b4ee, 32'h42bd73a4, 32'hc28bde81, 32'hc18d093e, 32'hc20b0137};
test_label[2867] = '{32'hc20b0137};
test_output[2867] = '{32'h43017a20};
/*############ DEBUG ############
test_input[22936:22943] = '{-74.5145000745, 43.30878281, -52.2692514296, 54.176687894, 94.7258616347, -69.934576719, -17.62951288, -34.751187025};
test_label[2867] = '{-34.751187025};
test_output[2867] = '{129.47704866};
############ END DEBUG ############*/
test_input[22944:22951] = '{32'h429862f4, 32'hc2b8c47e, 32'hc209d943, 32'hc1bd952c, 32'h428a9546, 32'h4186a8a0, 32'hc28b8ed0, 32'h40cc7e90};
test_label[2868] = '{32'h4186a8a0};
test_output[2868] = '{32'h426d729f};
/*############ DEBUG ############
test_input[22944:22951] = '{76.1932680931, -92.3837729487, -34.4621707751, -23.6978380446, 69.291548579, 16.832337379, -69.7789316654, 6.3904496918};
test_label[2868] = '{16.832337379};
test_output[2868] = '{59.3619362624};
############ END DEBUG ############*/
test_input[22952:22959] = '{32'h42bab6b5, 32'h42a13ce6, 32'h42911a1c, 32'hc2c1ca3e, 32'h42b2d0fc, 32'hc2506a1b, 32'h417df191, 32'h42a93ba2};
test_label[2869] = '{32'h42911a1c};
test_output[2869] = '{32'h41a699d3};
/*############ DEBUG ############
test_input[22952:22959] = '{93.3568499982, 80.6189453868, 72.550997929, -96.895003658, 89.4081742158, -52.1036170702, 15.8714764017, 84.6164720355};
test_label[2869] = '{72.550997929};
test_output[2869] = '{20.8251086142};
############ END DEBUG ############*/
test_input[22960:22967] = '{32'h400d25a4, 32'hc22137c6, 32'h42046087, 32'hc2aa1816, 32'hc2849a4a, 32'h4221aaac, 32'hc2bbc400, 32'h42b347cd};
test_label[2870] = '{32'hc22137c6};
test_output[2870] = '{32'h4301f1d8};
/*############ DEBUG ############
test_input[22960:22967] = '{2.20542228614, -40.3044678014, 33.0942660436, -85.0470412728, -66.3013479841, 40.4166712677, -93.8828087478, 89.6402382227};
test_label[2870] = '{-40.3044678014};
test_output[2870] = '{129.944706024};
############ END DEBUG ############*/
test_input[22968:22975] = '{32'h41d5432e, 32'h41de934e, 32'hc282106d, 32'h41eba1ca, 32'h4095d3a4, 32'h429d28ad, 32'hc2339eaf, 32'h41683860};
test_label[2871] = '{32'h4095d3a4};
test_output[2871] = '{32'h4293cb73};
/*############ DEBUG ############
test_input[22968:22975] = '{26.6578035342, 27.8219260344, -65.03208527, 29.4539987898, 4.68208487179, 78.5794429555, -44.9049630901, 14.5137631644};
test_label[2871] = '{4.68208487179};
test_output[2871] = '{73.8973580837};
############ END DEBUG ############*/
test_input[22976:22983] = '{32'h429731e7, 32'h410452ae, 32'hc2538a2d, 32'h42b1cfc3, 32'hc1b70a58, 32'h42c097b8, 32'h42924494, 32'h4201ac0b};
test_label[2872] = '{32'h4201ac0b};
test_output[2872] = '{32'h427f8407};
/*############ DEBUG ############
test_input[22976:22983] = '{75.5974636478, 8.27018585205, -52.8849389138, 88.9057865362, -22.880051139, 96.2963256132, 73.1339380824, 32.4180101289};
test_label[2872] = '{32.4180101289};
test_output[2872] = '{63.8789323584};
############ END DEBUG ############*/
test_input[22984:22991] = '{32'hc28d7721, 32'h42641e7f, 32'hc2823d6c, 32'h40d53627, 32'hc29af781, 32'hc2a31617, 32'hc20500df, 32'hc1f50b19};
test_label[2873] = '{32'h40d53627};
test_output[2873] = '{32'h424977ba};
/*############ DEBUG ############
test_input[22984:22991] = '{-70.7326770692, 57.0297824718, -65.1199628743, 6.66286037873, -77.4834079707, -81.5431474983, -33.2508503205, -30.6304189455};
test_label[2873] = '{6.66286037873};
test_output[2873] = '{50.3669220931};
############ END DEBUG ############*/
test_input[22992:22999] = '{32'h40f478e8, 32'h42930f33, 32'hc229b526, 32'hc262b083, 32'h3f87eb04, 32'hc09b9638, 32'h42029f68, 32'h425c393b};
test_label[2874] = '{32'hc229b526};
test_output[2874] = '{32'h42e7e9c7};
/*############ DEBUG ############
test_input[22992:22999] = '{7.6397591015, 73.5296896619, -42.4269034605, -56.672375163, 1.06185960231, -4.86208712879, 32.6556683161, 55.0558902875};
test_label[2874] = '{-42.4269034605};
test_output[2874] = '{115.956593132};
############ END DEBUG ############*/
test_input[23000:23007] = '{32'h41c5285b, 32'hc1f1eeca, 32'h4259988d, 32'hc2afe8bf, 32'hc205ce44, 32'h42b19457, 32'hc219c5f7, 32'h410bbaf2};
test_label[2875] = '{32'h42b19457};
test_output[2875] = '{32'h26b00000};
/*############ DEBUG ############
test_input[23000:23007] = '{24.6447048156, -30.2415955943, 54.3989738156, -87.9545853265, -33.4514329453, 88.7897230166, -38.4433246414, 8.73314133332};
test_label[2875] = '{88.7897230166};
test_output[2875] = '{1.22124532709e-15};
############ END DEBUG ############*/
test_input[23008:23015] = '{32'h408154f7, 32'hc09e945a, 32'h40d08662, 32'hc228b8d0, 32'hc1c199ac, 32'hc2b365ec, 32'hc1d45e11, 32'h422d368e};
test_label[2876] = '{32'hc2b365ec};
test_output[2876] = '{32'h4305009a};
/*############ DEBUG ############
test_input[23008:23015] = '{4.04162171896, -4.95560933114, 6.5164039202, -42.1804813996, -24.2000347529, -89.6990693046, -26.5459312848, 43.3032756579};
test_label[2876] = '{-89.6990693046};
test_output[2876] = '{133.002344963};
############ END DEBUG ############*/
test_input[23016:23023] = '{32'h4185a305, 32'h41add87c, 32'h429b2681, 32'h429485b9, 32'h42bb3cfe, 32'hc2b47ae6, 32'hc275cc40, 32'hc2aacfe7};
test_label[2877] = '{32'h4185a305};
test_output[2877] = '{32'h4299d43d};
/*############ DEBUG ############
test_input[23016:23023] = '{16.7045992814, 21.7307055096, 77.5752009608, 74.2611799872, 93.619123334, -90.2400346724, -61.4494628343, -85.4060564035};
test_label[2877] = '{16.7045992814};
test_output[2877] = '{76.9145241642};
############ END DEBUG ############*/
test_input[23024:23031] = '{32'hc2872a14, 32'h41102ca9, 32'hc267af90, 32'h422104e0, 32'h4255b650, 32'hc296d85c, 32'h42b1f86c, 32'h41e3f076};
test_label[2878] = '{32'h4255b650};
test_output[2878] = '{32'h420e3a88};
/*############ DEBUG ############
test_input[23024:23031] = '{-67.5821842588, 9.01090314331, -57.921449159, 40.2547604737, 53.4280385762, -75.4225732435, 88.9851994954, 28.4924116942};
test_label[2878] = '{53.4280385762};
test_output[2878] = '{35.5571609192};
############ END DEBUG ############*/
test_input[23032:23039] = '{32'h4290c64e, 32'h4242a333, 32'h409a3529, 32'hc27da860, 32'h421ecde1, 32'h4154bc57, 32'hc2982391, 32'hc1ac37ae};
test_label[2879] = '{32'h4154bc57};
test_output[2879] = '{32'h426c5d87};
/*############ DEBUG ############
test_input[23032:23039] = '{72.387315267, 48.6593754047, 4.81898943692, -63.4144275036, 39.7010540435, 13.2959809571, -76.0694669153, -21.5271875655};
test_label[2879] = '{13.2959809571};
test_output[2879] = '{59.09133431};
############ END DEBUG ############*/
test_input[23040:23047] = '{32'h422e288c, 32'h418dddf1, 32'h42893908, 32'h424b758a, 32'h42760f53, 32'hc295d610, 32'h419b999a, 32'hc2b4d11b};
test_label[2880] = '{32'hc295d610};
test_output[2880] = '{32'h430f87c2};
/*############ DEBUG ############
test_input[23040:23047] = '{43.5395976558, 17.7333695509, 68.6113857607, 50.8647850879, 61.5149641878, -74.91808895, 19.4500010139, -90.4084086065};
test_label[2880] = '{-74.91808895};
test_output[2880] = '{143.53030245};
############ END DEBUG ############*/
test_input[23048:23055] = '{32'h42bae2b0, 32'hc11e3691, 32'hc285a210, 32'h41f5ff1c, 32'hc258794b, 32'h426b7273, 32'h41f039e9, 32'h41b048bc};
test_label[2881] = '{32'hc285a210};
test_output[2881] = '{32'h43204260};
/*############ DEBUG ############
test_input[23048:23055] = '{93.4427471366, -9.88832155819, -66.8165303106, 30.7495648232, -54.1184489315, 58.8617651566, 30.0282770109, 22.0355151183};
test_label[2881] = '{-66.8165303106};
test_output[2881] = '{160.259277447};
############ END DEBUG ############*/
test_input[23056:23063] = '{32'h41e41e39, 32'hc203e5cf, 32'hc03ff771, 32'h40d53096, 32'hc2ac4f0d, 32'hc1cb59ae, 32'hc2a34e1e, 32'hc2ab615d};
test_label[2882] = '{32'hc03ff771};
test_output[2882] = '{32'h41fc1d28};
/*############ DEBUG ############
test_input[23056:23063] = '{28.514757893, -32.9744228208, -2.99947764383, 6.66218081806, -86.1543954932, -25.4187896905, -81.6525740187, -85.6901641491};
test_label[2882] = '{-2.99947764383};
test_output[2882] = '{31.5142355372};
############ END DEBUG ############*/
test_input[23064:23071] = '{32'hc16e1087, 32'h42a0c058, 32'hc2ba4afa, 32'hc279c2c5, 32'hc03c54b7, 32'h427ea38a, 32'hc22636d2, 32'h42a2d8cc};
test_label[2883] = '{32'hc22636d2};
test_output[2883] = '{32'h42f68e22};
/*############ DEBUG ############
test_input[23064:23071] = '{-14.8790350265, 80.3756740598, -93.1464355646, -62.4402027425, -2.94267048354, 63.659706143, -41.5535338076, 81.4234318292};
test_label[2883] = '{-41.5535338076};
test_output[2883] = '{123.277605856};
############ END DEBUG ############*/
test_input[23072:23079] = '{32'hc2751e46, 32'hc26e7233, 32'h42855de7, 32'h428b7517, 32'hbf7ea94c, 32'h426bf694, 32'h421f737f, 32'h42ad2fce};
test_label[2884] = '{32'h42ad2fce};
test_output[2884] = '{32'h33554438};
/*############ DEBUG ############
test_input[23072:23079] = '{-61.2795647143, -59.611521584, 66.6834003882, 69.7286939978, -0.994770766069, 58.990797198, 39.8627898026, 86.5933669905};
test_label[2884] = '{86.5933669905};
test_output[2884] = '{4.96549714795e-08};
############ END DEBUG ############*/
test_input[23080:23087] = '{32'h4226a3c1, 32'h416e89cb, 32'hc253f546, 32'h42b89474, 32'hc248f0dd, 32'hc29bd3a8, 32'h42bfe10b, 32'h408692ef};
test_label[2885] = '{32'h42b89474};
test_output[2885] = '{32'h406b3782};
/*############ DEBUG ############
test_input[23080:23087] = '{41.6599176415, 14.9086407324, -52.9895250362, 92.2899440057, -50.2352198339, -77.9133935781, 95.9395375253, 4.20543611739};
test_label[2885] = '{92.2899440057};
test_output[2885] = '{3.67526291925};
############ END DEBUG ############*/
test_input[23088:23095] = '{32'h4296aa25, 32'h42bd041d, 32'h41ca2319, 32'h42994d62, 32'h427a069d, 32'h42bd571d, 32'hc2899adf, 32'hc2bc6ae8};
test_label[2886] = '{32'h41ca2319};
test_output[2886] = '{32'h428c0969};
/*############ DEBUG ############
test_input[23088:23095] = '{75.3323167176, 94.508031073, 25.2671384674, 76.6511402781, 62.5064576835, 94.6701431137, -68.8024788907, -94.2087988043};
test_label[2886] = '{25.2671384674};
test_output[2886] = '{70.0183772651};
############ END DEBUG ############*/
test_input[23096:23103] = '{32'h4211fb24, 32'h42a01590, 32'h4219f854, 32'hc2b8e329, 32'hc2ae160e, 32'hc29c63cf, 32'h421ec6e9, 32'h42247fd4};
test_label[2887] = '{32'hc2b8e329};
test_output[2887] = '{32'h432c7c5d};
/*############ DEBUG ############
test_input[23096:23103] = '{36.4952552967, 80.0421159443, 38.4925084193, -92.443675178, -87.043077874, -78.1949407383, 39.6942482626, 41.1248312409};
test_label[2887] = '{-92.443675178};
test_output[2887] = '{172.485791122};
############ END DEBUG ############*/
test_input[23104:23111] = '{32'h40fe6053, 32'hc2c39170, 32'h412fdb26, 32'hc276be3a, 32'h4189f7d7, 32'hc05f0471, 32'h42b187d7, 32'h428adaab};
test_label[2888] = '{32'h4189f7d7};
test_output[2888] = '{32'h428f09e1};
/*############ DEBUG ############
test_input[23104:23111] = '{7.94925827986, -97.7840605858, 10.9910034997, -61.6857685879, 17.2460153807, -3.4846461214, 88.7653128274, 69.4270870987};
test_label[2888] = '{17.2460153807};
test_output[2888] = '{71.5192974507};
############ END DEBUG ############*/
test_input[23112:23119] = '{32'hc17ee150, 32'hc1894c72, 32'h40a1a3ca, 32'hbfae128f, 32'hc23235a8, 32'h4264c592, 32'hc279fdfb, 32'hc200dcbb};
test_label[2889] = '{32'hc23235a8};
test_output[2889] = '{32'h42cb7d9d};
/*############ DEBUG ############
test_input[23112:23119] = '{-15.9300082124, -17.1623261457, 5.05124398755, -1.35994130405, -44.5523968044, 57.1929384354, -62.498027477, -32.2155562039};
test_label[2889] = '{-44.5523968044};
test_output[2889] = '{101.74533524};
############ END DEBUG ############*/
test_input[23120:23127] = '{32'hc2126ca7, 32'h426c9bf3, 32'hc118eb1f, 32'hc1e27ead, 32'hc261886d, 32'h42c0d851, 32'h4292014e, 32'hc0ce52fd};
test_label[2890] = '{32'h426c9bf3};
test_output[2890] = '{32'h421514af};
/*############ DEBUG ############
test_input[23120:23127] = '{-36.6061071361, 59.1522927013, -9.55740239543, -28.3118543081, -56.3832266292, 96.4224922374, 73.0025510231, -6.44763021206};
test_label[2890] = '{59.1522927013};
test_output[2890] = '{37.2701995362};
############ END DEBUG ############*/
test_input[23128:23135] = '{32'h41e2ad6c, 32'h42b4dae6, 32'hc18d1301, 32'hc24900b2, 32'h41856893, 32'h424bc890, 32'hc29b20bb, 32'hc18317b5};
test_label[2891] = '{32'h424bc890};
test_output[2891] = '{32'h421ded3d};
/*############ DEBUG ############
test_input[23128:23135] = '{28.3346789247, 90.4275388367, -17.634279632, -50.2506785939, 16.6760606823, 50.9458602043, -77.5639295592, -16.3865757371};
test_label[2891] = '{50.9458602043};
test_output[2891] = '{39.4816786324};
############ END DEBUG ############*/
test_input[23136:23143] = '{32'h42783ffb, 32'hc20c79ec, 32'h410134eb, 32'hc288d430, 32'hc2a54604, 32'hc26cef5c, 32'h42b6d3db, 32'h421789b8};
test_label[2892] = '{32'h421789b8};
test_output[2892] = '{32'h42561dfe};
/*############ DEBUG ############
test_input[23136:23143] = '{62.0624796266, -35.1190633237, 8.07541943787, -68.4144306836, -82.6367467754, -59.2337493557, 91.4137799901, 37.8844894489};
test_label[2892] = '{37.8844894489};
test_output[2892] = '{53.5292905411};
############ END DEBUG ############*/
test_input[23144:23151] = '{32'h42939488, 32'hc2865762, 32'h42c0ba4a, 32'hc280e032, 32'h42a2a83b, 32'hc27fea23, 32'h428b6fd5, 32'h42a2f02a};
test_label[2893] = '{32'h42939488};
test_output[2893] = '{32'h41b4970a};
/*############ DEBUG ############
test_input[23144:23151] = '{73.7901001111, -67.1706715956, 96.3638494118, -64.4378841502, 81.3285769334, -63.9786473847, 69.7184239997, 81.4690699699};
test_label[2893] = '{73.7901001111};
test_output[2893] = '{22.573749936};
############ END DEBUG ############*/
test_input[23152:23159] = '{32'hc2b61c3b, 32'hc1e0ee51, 32'hc2855d75, 32'hc13a0757, 32'hc28715e6, 32'hc2c219b6, 32'h42ae41ca, 32'hc2a60f0d};
test_label[2894] = '{32'hc2855d75};
test_output[2894] = '{32'h4319cf9f};
/*############ DEBUG ############
test_input[23152:23159] = '{-91.0551403637, -28.1163652778, -66.6825315514, -11.6267920851, -67.5427722772, -97.0502178857, 87.1284933549, -83.0293945336};
test_label[2894] = '{-66.6825315514};
test_output[2894] = '{153.811024906};
############ END DEBUG ############*/
test_input[23160:23167] = '{32'h42a877ad, 32'h42125687, 32'hc247b524, 32'h41615f60, 32'h4284538d, 32'h42399e6e, 32'h42363ab8, 32'hc2818b31};
test_label[2895] = '{32'h42a877ad};
test_output[2895] = '{32'h3273d2c0};
/*############ DEBUG ############
test_input[23160:23167] = '{84.2337448534, 36.5844983009, -49.9268958367, 14.0857852189, 66.1631842637, 46.4047163287, 45.5573432393, -64.7718561416};
test_label[2895] = '{84.2337448534};
test_output[2895] = '{1.41923805938e-08};
############ END DEBUG ############*/
test_input[23168:23175] = '{32'hc2c0fcbf, 32'h42803c68, 32'h412a6d95, 32'hc125d507, 32'hc2606f2d, 32'h42c5470c, 32'h42c00935, 32'h4270fe9c};
test_label[2896] = '{32'h42c5470c};
test_output[2896] = '{32'h3d8fd080};
/*############ DEBUG ############
test_input[23168:23175] = '{-96.493648187, 64.1179780682, 10.6517534052, -10.3645088842, -56.1085688915, 98.638763603, 96.0179849968, 60.2486412101};
test_label[2896] = '{98.638763603};
test_output[2896] = '{0.0702219027023};
############ END DEBUG ############*/
test_input[23176:23183] = '{32'hc295dd2f, 32'h4092cee5, 32'hc232d3a7, 32'h429d0e17, 32'h429f2488, 32'hc2b4e498, 32'h4283aacb, 32'hc0135d29};
test_label[2897] = '{32'hc295dd2f};
test_output[2897] = '{32'h431ace15};
/*############ DEBUG ############
test_input[23176:23183] = '{-74.9319982233, 4.58775569781, -44.7066914388, 78.5275177345, 79.571347053, -90.4464757184, 65.8335835303, -2.30256100287};
test_label[2897] = '{-74.9319982233};
test_output[2897] = '{154.80500781};
############ END DEBUG ############*/
test_input[23184:23191] = '{32'hc227f534, 32'h4273fd3f, 32'hc276b977, 32'hc2c5d40a, 32'hc1e1883c, 32'hc1f097ea, 32'h41a64f3d, 32'hc2ad2bd0};
test_label[2898] = '{32'hc2c5d40a};
test_output[2898] = '{32'h431fe955};
/*############ DEBUG ############
test_input[23184:23191] = '{-41.9894550397, 60.9973101158, -61.6811194013, -98.914140888, -28.1915211065, -30.074176654, 20.7886909726, -86.5855708952};
test_label[2898] = '{-98.914140888};
test_output[2898] = '{159.911451004};
############ END DEBUG ############*/
test_input[23192:23199] = '{32'h426a50df, 32'hc1e55094, 32'h40f5a441, 32'h41455fc2, 32'h41c38f1e, 32'h42bb86e6, 32'h42a41148, 32'h3f342ab2};
test_label[2899] = '{32'h40f5a441};
test_output[2899] = '{32'h42ac2ca3};
/*############ DEBUG ############
test_input[23192:23199] = '{58.5789773107, -28.6643447202, 7.67630057992, 12.3358784974, 24.4448809409, 93.7634752097, 82.0337545723, 0.703776505736};
test_label[2899] = '{7.67630057992};
test_output[2899] = '{86.0871826807};
############ END DEBUG ############*/
test_input[23200:23207] = '{32'h42af3176, 32'h42a36e8d, 32'hc1d55e3e, 32'h42c510b8, 32'h41f8eb35, 32'h4236b8a2, 32'hc25f0a86, 32'h42c66709};
test_label[2900] = '{32'h42c510b8};
test_output[2900] = '{32'h3f8a8932};
/*############ DEBUG ############
test_input[23200:23207] = '{87.5966031919, 81.7159167349, -26.6710158574, 98.532657311, 31.1148479408, 45.6803042125, -55.7602779138, 99.2012439502};
test_label[2900] = '{98.532657311};
test_output[2900] = '{1.08231184989};
############ END DEBUG ############*/
test_input[23208:23215] = '{32'h4213c3f6, 32'hc2085af2, 32'hc2891a92, 32'hc2365c58, 32'hc1c83ed3, 32'hc27d24f4, 32'hc2c3036a, 32'h42c3ab2d};
test_label[2901] = '{32'h42c3ab2d};
test_output[2901] = '{32'h80000000};
/*############ DEBUG ############
test_input[23208:23215] = '{36.9413666017, -34.0888128731, -68.5518988182, -45.5901783927, -25.0306764628, -63.2860855532, -97.5066701307, 97.8343258321};
test_label[2901] = '{97.8343258321};
test_output[2901] = '{-0.0};
############ END DEBUG ############*/
test_input[23216:23223] = '{32'hc242d03b, 32'h4170df8a, 32'h42ad7704, 32'hc19b9d24, 32'h4291ac3d, 32'hbf81795b, 32'h42a3e2a1, 32'h42454ba3};
test_label[2902] = '{32'h4291ac3d};
test_output[2902] = '{32'h415e7822};
/*############ DEBUG ############
test_input[23216:23223] = '{-48.7033499053, 15.0545746351, 86.7324491654, -19.4517290769, 72.8364008, -1.01151598091, 81.9426350218, 49.3238636149};
test_label[2902] = '{72.8364008};
test_output[2902] = '{13.9043289119};
############ END DEBUG ############*/
test_input[23224:23231] = '{32'h4270626e, 32'hc1f83d6d, 32'h426f86da, 32'h42adf551, 32'h429c00c2, 32'hc2a8d2ca, 32'h4127d7cd, 32'h42448894};
test_label[2903] = '{32'h4270626e};
test_output[2903] = '{32'h41d710aa};
/*############ DEBUG ############
test_input[23224:23231] = '{60.0961239868, -31.0299935235, 59.8816924713, 86.9791347028, 78.0014785015, -84.4116954953, 10.4901860344, 49.1333777112};
test_label[2903] = '{60.0961239868};
test_output[2903] = '{26.8831369063};
############ END DEBUG ############*/
test_input[23232:23239] = '{32'hc25d2981, 32'hc2a1c77f, 32'h42ae5cb6, 32'hc1936020, 32'h42a4ab5d, 32'hc2baa83d, 32'hc1c69b10, 32'hc2a75e27};
test_label[2904] = '{32'hc2baa83d};
test_output[2904] = '{32'h4334847a};
/*############ DEBUG ############
test_input[23232:23239] = '{-55.2905323732, -80.8896377156, 87.1810791397, -18.421936891, 82.3346916879, -93.3285868012, -24.825714299, -83.6838937311};
test_label[2904] = '{-93.3285868012};
test_output[2904] = '{180.517491947};
############ END DEBUG ############*/
test_input[23240:23247] = '{32'h418d9a1f, 32'hc267265e, 32'h42960fb9, 32'hc291a525, 32'hc2a23292, 32'hc2950961, 32'hc25d4749, 32'h42bcd7f2};
test_label[2905] = '{32'hc2a23292};
test_output[2905] = '{32'h432f8542};
/*############ DEBUG ############
test_input[23240:23247] = '{17.7002551706, -57.7874694112, 75.0307104886, -72.8225451692, -81.0987710633, -74.5183163645, -55.3196141672, 94.4217675288};
test_label[2905] = '{-81.0987710633};
test_output[2905] = '{175.520538596};
############ END DEBUG ############*/
test_input[23248:23255] = '{32'hc29a2eca, 32'h42bd0567, 32'hc2a50579, 32'h42c11dda, 32'hc214a303, 32'h42c6e6de, 32'h42938111, 32'h426e866d};
test_label[2906] = '{32'hc214a303};
test_output[2906] = '{32'h4308abba};
/*############ DEBUG ############
test_input[23248:23255] = '{-77.0913846867, 94.5105530998, -82.5106910226, 96.5583045566, -37.1591900808, 99.4509113658, 73.7520845546, 59.6312770228};
test_label[2906] = '{-37.1591900808};
test_output[2906] = '{136.67080471};
############ END DEBUG ############*/
test_input[23256:23263] = '{32'hc2883ff8, 32'h424d9e70, 32'h428ba23e, 32'hc1f4614b, 32'hc1fa14ae, 32'h40bc216d, 32'h429a06d4, 32'hc28de308};
test_label[2907] = '{32'hc1f4614b};
test_output[2907] = '{32'h42d71f89};
/*############ DEBUG ############
test_input[23256:23263] = '{-68.1249402958, 51.4047243848, 69.8168814891, -30.5475069592, -31.2600983643, 5.87908030964, 77.0133389738, -70.9434182577};
test_label[2907] = '{-30.5475069592};
test_output[2907] = '{107.561594888};
############ END DEBUG ############*/
test_input[23264:23271] = '{32'h428f52e7, 32'h42a35455, 32'hc29c032a, 32'hc285642c, 32'hc2530c32, 32'hc211ce1c, 32'h4209ea09, 32'h42aa35aa};
test_label[2908] = '{32'h428f52e7};
test_output[2908] = '{32'h4157975a};
/*############ DEBUG ############
test_input[23264:23271] = '{71.6619181617, 81.6647129212, -78.0061832689, -66.69565179, -52.7619080366, -36.451279754, 34.4785509786, 85.1048092899};
test_label[2908] = '{71.6619181617};
test_output[2908] = '{13.4744508854};
############ END DEBUG ############*/
test_input[23272:23279] = '{32'h4296f430, 32'h41662575, 32'h4204e81d, 32'h4198164b, 32'hc29ca458, 32'h425e5c1c, 32'h41c3d920, 32'h423093b9};
test_label[2909] = '{32'h4296f430};
test_output[2909] = '{32'h311e975e};
/*############ DEBUG ############
test_input[23272:23279] = '{75.476929272, 14.3841444497, 33.2266714924, 19.0108845432, -78.3209871966, 55.5899503603, 24.4810178383, 44.1442589089};
test_label[2909] = '{75.476929272};
test_output[2909] = '{2.30780672616e-09};
############ END DEBUG ############*/
test_input[23280:23287] = '{32'h42747175, 32'hc159e350, 32'hc2c51597, 32'hc21e442c, 32'h4239bdd6, 32'hc18e77ff, 32'hc290ef31, 32'h418d30b0};
test_label[2910] = '{32'hc2c51597};
test_output[2910] = '{32'h431fa729};
/*############ DEBUG ############
test_input[23280:23287] = '{61.1107982164, -13.6179963718, -98.5421686325, -39.56657517, 46.4353875125, -17.8085909694, -72.467172659, 17.6487730059};
test_label[2910] = '{-98.5421686325};
test_output[2910] = '{159.652967272};
############ END DEBUG ############*/
test_input[23288:23295] = '{32'hc2c601b6, 32'h42976608, 32'h4281a5c1, 32'hc2b2c324, 32'h4283cf38, 32'hc1ec1533, 32'h428b0996, 32'hc24b2209};
test_label[2911] = '{32'h42976608};
test_output[2911] = '{32'h3b0c5b05};
/*############ DEBUG ############
test_input[23288:23295] = '{-99.0033443402, 75.6992796619, 64.8237418622, -89.3811375663, 65.9047216951, -29.5103512353, 69.5187255973, -50.7832392786};
test_label[2911] = '{75.6992796619};
test_output[2911] = '{0.00214165556172};
############ END DEBUG ############*/
test_input[23296:23303] = '{32'hc2b90e20, 32'hc294a4ae, 32'hc07d9f8e, 32'hc2a9c35d, 32'h42a19337, 32'h421c9c0f, 32'hc283bed1, 32'h41ae5162};
test_label[2912] = '{32'hc07d9f8e};
test_output[2912] = '{32'h42a98033};
/*############ DEBUG ############
test_input[23296:23303] = '{-92.5275880528, -74.321637263, -3.96286337614, -84.8815688681, 80.7875290812, 39.1523992086, -65.8726904829, 21.7897372104};
test_label[2912] = '{-3.96286337614};
test_output[2912] = '{84.7503924574};
############ END DEBUG ############*/
test_input[23304:23311] = '{32'hc13fee23, 32'hc2c7f0b9, 32'h422bb8c5, 32'hc2216383, 32'hc205aa3e, 32'hc28fc149, 32'h4199d31f, 32'hc22d3adf};
test_label[2913] = '{32'hc28fc149};
test_output[2913] = '{32'h42e59dac};
/*############ DEBUG ############
test_input[23304:23311] = '{-11.9956388544, -99.9701591077, 42.9304402315, -40.3471793427, -33.4162536076, -71.8775108559, 19.2280869456, -43.3074922704};
test_label[2913] = '{-71.8775108559};
test_output[2913] = '{114.807951087};
############ END DEBUG ############*/
test_input[23312:23319] = '{32'hc27b4f9a, 32'h42917d99, 32'hc040cfcb, 32'h426a48f4, 32'hc21059ad, 32'h429dccf1, 32'h42bf26de, 32'h42c141a9};
test_label[2914] = '{32'hc040cfcb};
test_output[2914] = '{32'h42c7e17a};
/*############ DEBUG ############
test_input[23312:23319] = '{-62.8277342042, 72.7453099398, -3.01268274339, 58.5712416985, -36.0875739453, 78.9002785455, 95.5759117012, 96.6282438157};
test_label[2914] = '{-3.01268274339};
test_output[2914] = '{99.940381033};
############ END DEBUG ############*/
test_input[23320:23327] = '{32'hc2819f32, 32'hc0a0995e, 32'h421df164, 32'h41933cff, 32'hc2b2e562, 32'hc2bf89a3, 32'h41a42822, 32'h4217a24d};
test_label[2915] = '{32'h421df164};
test_output[2915] = '{32'h3e40446c};
/*############ DEBUG ############
test_input[23320:23327] = '{-64.8109312329, -5.0187215545, 39.4857337221, 18.4047825141, -89.4480123065, -95.7688212463, 20.5195961415, 37.9084973013};
test_label[2915] = '{39.4857337221};
test_output[2915] = '{0.187761003217};
############ END DEBUG ############*/
test_input[23328:23335] = '{32'h42b07c17, 32'hc295d0be, 32'hc1c74875, 32'hc19f1c78, 32'h42a8483e, 32'hc2b23743, 32'hc28e8f99, 32'hc2c679b1};
test_label[2916] = '{32'hc2b23743};
test_output[2916] = '{32'h43315de1};
/*############ DEBUG ############
test_input[23328:23335] = '{88.242363353, -74.9077018118, -24.910378746, -19.8889012006, 84.1410974848, -89.107930062, -71.2804670743, -99.2376818213};
test_label[2916] = '{-89.107930062};
test_output[2916] = '{177.366709638};
############ END DEBUG ############*/
test_input[23336:23343] = '{32'hc278a830, 32'h42a015d5, 32'h42c243db, 32'h42c54544, 32'h41957eb1, 32'h42b14dfd, 32'hc20b3c2b, 32'h42bd4e6e};
test_label[2917] = '{32'h42a015d5};
test_output[2917] = '{32'h41967849};
/*############ DEBUG ############
test_input[23336:23343] = '{-62.164244477, 80.0426369076, 97.1325340111, 98.635283956, 18.6868614342, 88.6523236109, -34.8087569751, 94.653183502};
test_label[2917] = '{80.0426369076};
test_output[2917] = '{18.8087337814};
############ END DEBUG ############*/
test_input[23344:23351] = '{32'hc1b8531f, 32'hc1f49b6d, 32'hc1019281, 32'h4210939a, 32'hc11b78c6, 32'hc2b2efe7, 32'hbfb769a4, 32'hc1b96acf};
test_label[2918] = '{32'hc11b78c6};
test_output[2918] = '{32'h423771cb};
/*############ DEBUG ############
test_input[23344:23351] = '{-23.0405859091, -30.5758912674, -8.09826779151, 36.1441410702, -9.71698555761, -89.4685569985, -1.43291145142, -23.1771523433};
test_label[2918] = '{-9.71698555761};
test_output[2918] = '{45.8611266278};
############ END DEBUG ############*/
test_input[23352:23359] = '{32'h42952991, 32'h427ed16f, 32'h40e3c9a2, 32'h42b79556, 32'h426597f6, 32'h42bef404, 32'hc22326a2, 32'h42888443};
test_label[2919] = '{32'h42b79556};
test_output[2919] = '{32'h406d6be1};
/*############ DEBUG ############
test_input[23352:23359] = '{74.5811875354, 63.7045255397, 7.11836336106, 91.791672453, 57.3983988752, 95.47659242, -40.787728977, 68.258320586};
test_label[2919] = '{91.791672453};
test_output[2919] = '{3.70970934002};
############ END DEBUG ############*/
test_input[23360:23367] = '{32'h42c7561f, 32'h42a576ce, 32'hc24a8cc4, 32'hc1b07d81, 32'hc2550f4c, 32'h42140998, 32'hc2b493b9, 32'h4261b1d6};
test_label[2920] = '{32'hc2b493b9};
test_output[2920] = '{32'h433df4ec};
/*############ DEBUG ############
test_input[23360:23367] = '{99.6682045458, 82.7320368468, -50.6374661708, -22.0612806156, -53.2649389794, 37.0093691305, -90.2885226962, 56.4236693883};
test_label[2920] = '{-90.2885226962};
test_output[2920] = '{189.956727286};
############ END DEBUG ############*/
test_input[23368:23375] = '{32'hc2a83b6b, 32'h42b72a3e, 32'hc1107a6c, 32'h42bf8348, 32'hc15c07e4, 32'hc2a17359, 32'h4056c78f, 32'hc1f1cbf6};
test_label[2921] = '{32'hc15c07e4};
test_output[2921] = '{32'h42db0c16};
/*############ DEBUG ############
test_input[23368:23375] = '{-84.1160490121, 91.5825058777, -9.02988772273, 95.7564060297, -13.7519261841, -80.7252902885, 3.35593016764, -30.2245908326};
test_label[2921] = '{-13.7519261841};
test_output[2921] = '{109.523607068};
############ END DEBUG ############*/
test_input[23376:23383] = '{32'h4227d031, 32'hc287536d, 32'hc26b1ea1, 32'hc2c2a9b8, 32'hc161bf79, 32'h42b65f42, 32'hc2bc7fb9, 32'hc241929e};
test_label[2922] = '{32'hc241929e};
test_output[2922] = '{32'h430b9449};
/*############ DEBUG ############
test_input[23376:23383] = '{41.9533109013, -67.6629411975, -58.7799119939, -97.3314787654, -14.1092457881, 91.1860520599, -94.2494557423, -48.3931801};
test_label[2922] = '{-48.3931801};
test_output[2922] = '{139.57923216};
############ END DEBUG ############*/
test_input[23384:23391] = '{32'hc2ba97e3, 32'hc1db22ac, 32'hc1397273, 32'hc29309be, 32'hc201313c, 32'hc2676e0c, 32'h42a74ad1, 32'hc28af7af};
test_label[2923] = '{32'hc28af7af};
test_output[2923] = '{32'h43192140};
/*############ DEBUG ############
test_input[23384:23391] = '{-93.2966514291, -27.3919299747, -11.59044123, -73.5190286366, -32.2980813706, -57.8574659978, 83.6461281065, -69.4837563138};
test_label[2923] = '{-69.4837563138};
test_output[2923] = '{153.12988442};
############ END DEBUG ############*/
test_input[23392:23399] = '{32'h41ea4e70, 32'h4275b4ec, 32'h426d4475, 32'h421ca9a5, 32'h428e75a0, 32'hc19449da, 32'hc28bf7cf, 32'hc274bd43};
test_label[2924] = '{32'h4275b4ec};
test_output[2924] = '{32'h411cd994};
/*############ DEBUG ############
test_input[23392:23399] = '{29.2882995854, 61.4266809055, 59.316852481, 39.1656688639, 71.2297389333, -18.5360594806, -69.9840039061, -61.1848245732};
test_label[2924] = '{61.4266809055};
test_output[2924] = '{9.80312001157};
############ END DEBUG ############*/
test_input[23400:23407] = '{32'hc2a38727, 32'h42a88da4, 32'hc25c1097, 32'h42b665b0, 32'h423311fa, 32'h42664e7e, 32'hc0dfe040, 32'h40240397};
test_label[2925] = '{32'h42664e7e};
test_output[2925] = '{32'h42067de5};
/*############ DEBUG ############
test_input[23400:23407] = '{-81.7639692153, 84.2766409402, -55.0162006871, 91.19860743, 44.7675558115, 57.5766507369, -6.9961241931, 2.56271920736};
test_label[2925] = '{57.5766507369};
test_output[2925] = '{33.6229420967};
############ END DEBUG ############*/
test_input[23408:23415] = '{32'hc29a2e15, 32'hc2bdbfc7, 32'h4275e9a7, 32'h426c35a1, 32'h41a9d7f0, 32'hc2b213c5, 32'h423c1933, 32'hc18f72cb};
test_label[2926] = '{32'hc29a2e15};
test_output[2926] = '{32'h430aa724};
/*############ DEBUG ############
test_input[23408:23415] = '{-77.0900042725, -94.8745655593, 61.4781755556, 59.052370115, 21.2304388762, -89.0386121722, 47.0246080507, -17.931050742};
test_label[2926] = '{-77.0900042725};
test_output[2926] = '{138.652895366};
############ END DEBUG ############*/
test_input[23416:23423] = '{32'h42bd5eed, 32'h42a3d473, 32'h42c18b7f, 32'h42aa194b, 32'h41a5a1c0, 32'hc2697acb, 32'hc0bfb98c, 32'hc17f3782};
test_label[2927] = '{32'h42a3d473};
test_output[2927] = '{32'h416f9766};
/*############ DEBUG ############
test_input[23416:23423] = '{94.6854023119, 81.9149389596, 96.7724537701, 85.0494023338, 20.7039788637, -58.3699139722, -5.9913999111, -15.9510520723};
test_label[2927] = '{81.9149389596};
test_output[2927] = '{14.9744626781};
############ END DEBUG ############*/
test_input[23424:23431] = '{32'hc29911b3, 32'h4280a48c, 32'h4288dc97, 32'hc20f6262, 32'hc25c73be, 32'h421f73c5, 32'hc210fd42, 32'h423e5db9};
test_label[2928] = '{32'h4280a48c};
test_output[2928] = '{32'h40840612};
/*############ DEBUG ############
test_input[23424:23431] = '{-76.5345677829, 64.3213807184, 68.4308384282, -35.8460765785, -55.1130300141, 39.8630546574, -36.2473206509, 47.591526053};
test_label[2928] = '{64.3213807184};
test_output[2928] = '{4.1257410887};
############ END DEBUG ############*/
test_input[23432:23439] = '{32'hc2ac484b, 32'h424c65f7, 32'h42a875c9, 32'hc0ad3016, 32'h42854302, 32'hc1a243ad, 32'hc279b9d7, 32'h4171c31c};
test_label[2929] = '{32'h4171c31c};
test_output[2929] = '{32'h428a3d66};
/*############ DEBUG ############
test_input[23432:23439] = '{-86.1411966635, 51.0995766264, 84.230051034, -5.41211965442, 66.6308725567, -20.2830455294, -62.4314831181, 15.1101337942};
test_label[2929] = '{15.1101337942};
test_output[2929] = '{69.1199172626};
############ END DEBUG ############*/
test_input[23440:23447] = '{32'h426e435f, 32'h42b90208, 32'hc20a8b82, 32'h429a80be, 32'h42bc0a2a, 32'h428da02d, 32'hc1d52dc9, 32'hc2be9c00};
test_label[2930] = '{32'hc2be9c00};
test_output[2930] = '{32'h433d85e8};
/*############ DEBUG ############
test_input[23440:23447] = '{59.5657928198, 92.5039640238, -34.6362393996, 77.2514468851, 94.0198534523, 70.8128451525, -26.6473568955, -95.3046840314};
test_label[2930] = '{-95.3046840314};
test_output[2930] = '{189.523070932};
############ END DEBUG ############*/
test_input[23448:23455] = '{32'hc2632222, 32'h4265e025, 32'hc0e875d8, 32'hc26978c5, 32'h4157ff4d, 32'h42763c69, 32'hc142d394, 32'hc290fd32};
test_label[2931] = '{32'hc142d394};
test_output[2931] = '{32'h42938127};
/*############ DEBUG ############
test_input[23448:23455] = '{-56.7833311332, 57.4688915353, -7.26438520048, -58.3679408574, 13.4998297015, 61.5589951438, -12.1766548662, -72.4945192418};
test_label[2931] = '{-12.1766548662};
test_output[2931] = '{73.752248981};
############ END DEBUG ############*/
test_input[23456:23463] = '{32'h4120be9f, 32'h421f6358, 32'h42adf7db, 32'hc28ef615, 32'h4274a05b, 32'h41852fb8, 32'h420e154c, 32'hc2498c62};
test_label[2932] = '{32'h4274a05b};
test_output[2932] = '{32'h41ce9eb6};
/*############ DEBUG ############
test_input[23456:23463] = '{10.0465380785, 39.8470166122, 86.9840913941, -71.4806265493, 61.1565956609, 16.6482997937, 35.5207970533, -50.3870927189};
test_label[2932] = '{61.1565956609};
test_output[2932] = '{25.8274957332};
############ END DEBUG ############*/
test_input[23464:23471] = '{32'hc21c7e2c, 32'hc1c71f4c, 32'h418ba987, 32'hc2223ba7, 32'h4225833c, 32'h425d84ba, 32'hc25a4f5c, 32'hc1929ec6};
test_label[2933] = '{32'hc1929ec6};
test_output[2933] = '{32'h42936a0f};
/*############ DEBUG ############
test_input[23464:23471] = '{-39.1232156533, -24.8902819621, 17.4577775333, -40.5582553849, 41.3781591679, 55.3796161132, -54.5774982229, -18.3275253965};
test_label[2933] = '{-18.3275253965};
test_output[2933] = '{73.70714234};
############ END DEBUG ############*/
test_input[23472:23479] = '{32'hc22fd671, 32'hc2b98964, 32'hc2bcff4b, 32'h40c579f8, 32'hc28df079, 32'hc28b4c7d, 32'hc24d3869, 32'h412e7a9b};
test_label[2934] = '{32'hc24d3869};
test_output[2934] = '{32'h4278e006};
/*############ DEBUG ############
test_input[23472:23479] = '{-43.9594144324, -92.7683441787, -94.4986183152, 6.17113858578, -70.9696727228, -69.6493893082, -51.3050862186, 10.9049333503};
test_label[2934] = '{-51.3050862186};
test_output[2934] = '{62.2187741754};
############ END DEBUG ############*/
test_input[23480:23487] = '{32'hc2c529d0, 32'h40d633ca, 32'h41e144ee, 32'h428c21c5, 32'h41e5a63f, 32'hc25c29c1, 32'h4253277b, 32'h42bf015a};
test_label[2935] = '{32'h42bf015a};
test_output[2935] = '{32'h2d1ddf80};
/*############ DEBUG ############
test_input[23480:23487] = '{-98.5816636883, 6.69382199173, 28.1586569601, 70.0659599274, 28.7061749551, -55.0407751664, 52.7885537074, 95.5026432338};
test_label[2935] = '{95.5026432338};
test_output[2935] = '{8.97404373039e-12};
############ END DEBUG ############*/
test_input[23488:23495] = '{32'hc268e725, 32'h42988865, 32'hc2783f77, 32'h4187ac06, 32'h429e6618, 32'h425eec95, 32'hc2b45898, 32'h411021c7};
test_label[2936] = '{32'h4187ac06};
test_output[2936] = '{32'h42792b4a};
/*############ DEBUG ############
test_input[23488:23495] = '{-58.2257281118, 76.2663918272, -62.0619759664, 16.9589951444, 79.1994004765, 55.7310376451, -90.1730343429, 9.00824642285};
test_label[2936] = '{16.9589951444};
test_output[2936] = '{62.2922732566};
############ END DEBUG ############*/
test_input[23496:23503] = '{32'hc2018267, 32'h42ba8bd6, 32'hc1bd5220, 32'h42bc0fc8, 32'hc29fe0b6, 32'hc27922a4, 32'hc2c0777e, 32'h4285bf5e};
test_label[2937] = '{32'hc2c0777e};
test_output[2937] = '{32'h433ea60b};
/*############ DEBUG ############
test_input[23496:23503] = '{-32.3773477938, 93.2731195015, -23.6650991535, 94.0308256963, -79.9388882097, -62.2838288853, -96.2333815416, 66.8737620086};
test_label[2937] = '{-96.2333815416};
test_output[2937] = '{190.648612396};
############ END DEBUG ############*/
test_input[23504:23511] = '{32'hc288d424, 32'h411aed53, 32'h416abae9, 32'hc0b3d98e, 32'hc298a0c7, 32'hc28910b3, 32'h42c7d585, 32'h429bcb74};
test_label[2938] = '{32'h429bcb74};
test_output[2938] = '{32'h41b02844};
/*############ DEBUG ############
test_input[23504:23511] = '{-68.4143363159, 9.68294039959, 14.6706319197, -5.62030683011, -76.3140220146, -68.5326120264, 99.9170295388, 77.8973689448};
test_label[2938] = '{77.8973689448};
test_output[2938] = '{22.0196605942};
############ END DEBUG ############*/
test_input[23512:23519] = '{32'h429838fd, 32'h421d8555, 32'hc22868e4, 32'hc1a3781e, 32'h423c9a1a, 32'hc2a16478, 32'hc2418fc9, 32'h42b4a7c3};
test_label[2939] = '{32'h42b4a7c3};
test_output[2939] = '{32'h3533c954};
/*############ DEBUG ############
test_input[23512:23519] = '{76.1113084728, 39.38020638, -42.1024308055, -20.4336504336, 47.1504908251, -80.6962296467, -48.390417037, 90.3276594727};
test_label[2939] = '{90.3276594727};
test_output[2939] = '{6.6975669335e-07};
############ END DEBUG ############*/
test_input[23520:23527] = '{32'hc10b01ae, 32'h42c4e95b, 32'h42832cf6, 32'h40151bdb, 32'hc2a4d582, 32'hc29b11ee, 32'h41c56bb7, 32'h423a5b9d};
test_label[2940] = '{32'h42832cf6};
test_output[2940] = '{32'h420378cc};
/*############ DEBUG ############
test_input[23520:23527] = '{-8.68791009963, 98.4557748235, 65.5878105254, 2.32982507709, -82.4170088047, -77.5350188129, 24.6775954079, 46.5894661508};
test_label[2940] = '{65.5878105254};
test_output[2940] = '{32.8679642982};
############ END DEBUG ############*/
test_input[23528:23535] = '{32'h4288750f, 32'h3fed8a2f, 32'h42569fd4, 32'h42aa77fa, 32'hc13337a0, 32'h42aa271e, 32'hc1ae41b9, 32'h428a9915};
test_label[2941] = '{32'h42aa77fa};
test_output[2941] = '{32'h3f1e0748};
/*############ DEBUG ############
test_input[23528:23535] = '{68.2286291512, 1.85577951709, 53.6560839377, 85.2343305032, -11.2010800819, 85.0764045333, -21.7820910202, 69.298988436};
test_label[2941] = '{85.2343305032};
test_output[2941] = '{0.617298624696};
############ END DEBUG ############*/
test_input[23536:23543] = '{32'hc22576fa, 32'h42aad309, 32'h4183ea24, 32'h41a9242c, 32'hc28e460d, 32'hc2295952, 32'h40d8f4b7, 32'h4203b9b1};
test_label[2942] = '{32'h41a9242c};
test_output[2942] = '{32'h428089fe};
/*############ DEBUG ############
test_input[23536:23543] = '{-41.3661866306, 85.4121747346, 16.4893263309, 21.1426619956, -71.1368181639, -42.3372270834, 6.77987248823, 32.9313402847};
test_label[2942] = '{21.1426619956};
test_output[2942] = '{64.269512739};
############ END DEBUG ############*/
test_input[23544:23551] = '{32'hc1b06b20, 32'h42791a8a, 32'hc1ee5031, 32'hc29d09bf, 32'h42b84ef5, 32'hc28b6bac, 32'h41e3cafd, 32'hc2a075a6};
test_label[2943] = '{32'h42b84ef5};
test_output[2943] = '{32'h29ee0000};
/*############ DEBUG ############
test_input[23544:23551] = '{-22.0523064794, 62.2759181409, -29.7891556375, -78.5190344488, 92.1542108536, -69.7102999384, 28.4741149401, -80.2297845541};
test_label[2943] = '{92.1542108536};
test_output[2943] = '{1.05693231944e-13};
############ END DEBUG ############*/
test_input[23552:23559] = '{32'hc2801aaf, 32'hc2aa8e68, 32'hc2457302, 32'h42bad999, 32'hc2b6e530, 32'h422b87eb, 32'hc2861e40, 32'hc2297106};
test_label[2944] = '{32'hc2b6e530};
test_output[2944] = '{32'h4338df64};
/*############ DEBUG ############
test_input[23552:23559] = '{-64.0521146364, -85.2781338807, -49.3623141268, 93.4249917992, -91.4476306456, 42.8827326651, -67.0590810154, -42.3603732912};
test_label[2944] = '{-91.4476306456};
test_output[2944] = '{184.872622445};
############ END DEBUG ############*/
test_input[23560:23567] = '{32'hc247f8a5, 32'hc243067f, 32'h42680363, 32'h41f208c5, 32'h4158e7cb, 32'hc2346f02, 32'hc297302a, 32'hc2b9ffdb};
test_label[2945] = '{32'h4158e7cb};
test_output[2945] = '{32'h4231c970};
/*############ DEBUG ############
test_input[23560:23567] = '{-49.9928167923, -48.7563443877, 58.0033072516, 30.254281645, 13.55659051, -45.1084058424, -75.5940724238, -92.9997187268};
test_label[2945] = '{13.55659051};
test_output[2945] = '{44.4467167416};
############ END DEBUG ############*/
test_input[23568:23575] = '{32'h42c40a2d, 32'hc1207684, 32'hc251ef3e, 32'h42a7cbbf, 32'h42929aa4, 32'h4198af9e, 32'h4289f8f2, 32'hc1765e62};
test_label[2946] = '{32'hc1765e62};
test_output[2946] = '{32'h42e2d5f9};
/*############ DEBUG ############
test_input[23568:23575] = '{98.0198732312, -10.0289341281, -52.4836333165, 83.8979423285, 73.3020288766, 19.0857500578, 68.9862199855, -15.3980428543};
test_label[2946] = '{-15.3980428543};
test_output[2946] = '{113.417916822};
############ END DEBUG ############*/
test_input[23576:23583] = '{32'hc18c082b, 32'h4296a281, 32'hc286d927, 32'h42676106, 32'h423b3f72, 32'h420da2e1, 32'h42909a72, 32'h42970a95};
test_label[2947] = '{32'hc286d927};
test_output[2947] = '{32'h430f9031};
/*############ DEBUG ############
test_input[23576:23583] = '{-17.503987375, 75.3173926466, -67.4241248429, 57.8447484498, 46.8119599482, 35.4090602441, 72.3016520697, 75.520670317};
test_label[2947] = '{-67.4241248429};
test_output[2947] = '{143.563243547};
############ END DEBUG ############*/
test_input[23584:23591] = '{32'hc2758918, 32'h42b0a3b8, 32'h418cf135, 32'hc2bd02ea, 32'hbec180c5, 32'h42a33eda, 32'h42a59340, 32'hc2205f31};
test_label[2948] = '{32'h42a59340};
test_output[2948] = '{32'h40b131ea};
/*############ DEBUG ############
test_input[23584:23591] = '{-61.3838797157, 88.3197605263, 17.6177777033, -94.5056922074, -0.377935570847, 81.6227537784, 82.7875959783, -40.0929621354};
test_label[2948] = '{82.7875959783};
test_output[2948] = '{5.53734313161};
############ END DEBUG ############*/
test_input[23592:23599] = '{32'hc2b80696, 32'h41adcda5, 32'hc00c9419, 32'hc186f0a2, 32'h41cc098a, 32'hc27a6587, 32'hc28f1967, 32'hc124f82c};
test_label[2949] = '{32'hc28f1967};
test_output[2949] = '{32'h42c22759};
/*############ DEBUG ############
test_input[23592:23599] = '{-92.0128623259, 21.7254133157, -2.19653914689, -16.8674973332, 25.5046584489, -62.5991471386, -71.5496107423, -10.3105892814};
test_label[2949] = '{-71.5496107423};
test_output[2949] = '{97.0768521908};
############ END DEBUG ############*/
test_input[23600:23607] = '{32'h40a0da0e, 32'h429a242b, 32'h4200c5b2, 32'hbfbe343a, 32'h42a89707, 32'h42a5aeef, 32'hc1ddb420, 32'h429738ab};
test_label[2950] = '{32'hbfbe343a};
test_output[2950] = '{32'h42abfbc9};
/*############ DEBUG ############
test_input[23600:23607] = '{5.02661783069, 77.0706428082, 32.1930634559, -1.48596880227, 84.2949737578, 82.8416643185, -27.7129507773, 75.6106798314};
test_label[2950] = '{-1.48596880227};
test_output[2950] = '{85.9917650279};
############ END DEBUG ############*/
test_input[23608:23615] = '{32'hc205e490, 32'h42a081bf, 32'h427cb93b, 32'hc1a82f44, 32'h423bf4bb, 32'hc28adf88, 32'h427cdc8f, 32'h3feced0f};
test_label[2951] = '{32'h427cdc8f};
test_output[2951] = '{32'h41884ddf};
/*############ DEBUG ############
test_input[23608:23615] = '{-33.4732045793, 80.2534120613, 63.1808892649, -21.0230792396, 46.9889938845, -69.4365808557, 63.2153889622, 1.85098441775};
test_label[2951] = '{63.2153889622};
test_output[2951] = '{17.0380231774};
############ END DEBUG ############*/
test_input[23616:23623] = '{32'hc1c3d3b5, 32'h42197d06, 32'h42971db7, 32'h4234c278, 32'h42ae5938, 32'hc1fed18e, 32'h4214af89, 32'h42b70654};
test_label[2952] = '{32'h42197d06};
test_output[2952] = '{32'h42549ceb};
/*############ DEBUG ############
test_input[23616:23623] = '{-24.4783721787, 38.3720948411, 75.5580387377, 45.1899091005, 87.1742585425, -31.8523217641, 37.1714229222, 91.5123591367};
test_label[2952] = '{38.3720948411};
test_output[2952] = '{53.1532411618};
############ END DEBUG ############*/
test_input[23624:23631] = '{32'h427d5906, 32'h424269ea, 32'h423e4c23, 32'hc1b8af8e, 32'h4249363e, 32'h425061b8, 32'hc255e56c, 32'h4291bc7b};
test_label[2953] = '{32'h4249363e};
test_output[2953] = '{32'h41b48595};
/*############ DEBUG ############
test_input[23624:23631] = '{63.3369379462, 48.60343082, 47.5743505055, -23.0857207387, 50.3029727476, 52.095430361, -53.4740443607, 72.8681258168};
test_label[2953] = '{50.3029727476};
test_output[2953] = '{22.5652256211};
############ END DEBUG ############*/
test_input[23632:23639] = '{32'hc25b636c, 32'hc24b385b, 32'hc2abd27a, 32'hc297c266, 32'h42696ccc, 32'h41becbb2, 32'h4172d88a, 32'hc2ae2694};
test_label[2954] = '{32'hc2ae2694};
test_output[2954] = '{32'h43116e7d};
/*############ DEBUG ############
test_input[23632:23639] = '{-54.8470901717, -50.805035651, -85.9110836179, -75.8796835704, 58.3562467428, 23.8494609238, 15.1778655069, -87.0753490966};
test_label[2954] = '{-87.0753490966};
test_output[2954] = '{145.431595839};
############ END DEBUG ############*/
test_input[23640:23647] = '{32'h42918bb3, 32'hc2a813dd, 32'hc20665a4, 32'h426918f7, 32'h42bd62f4, 32'h4134183b, 32'hc259e284, 32'hc27fb829};
test_label[2955] = '{32'hc27fb829};
test_output[2955] = '{32'h431e9f84};
/*############ DEBUG ############
test_input[23640:23647] = '{72.7728468257, -84.0387925459, -33.5992595175, 58.2743811456, 94.6932651756, 11.2559152654, -54.4712071156, -63.929842777};
test_label[2955] = '{-63.929842777};
test_output[2955] = '{158.623107953};
############ END DEBUG ############*/
test_input[23648:23655] = '{32'h4224a1c5, 32'hc28af096, 32'hc21bbadb, 32'h42ab4e69, 32'hbf19ab9f, 32'h42c5a7a4, 32'hc277a345, 32'hc19e6aa3};
test_label[2956] = '{32'hc21bbadb};
test_output[2956] = '{32'h4309c289};
/*############ DEBUG ############
test_input[23648:23655] = '{41.1579791429, -69.4698906124, -38.9324748333, 85.6531435758, -0.600274959737, 98.8274227228, -61.9094432612, -19.8020682114};
test_label[2956] = '{-38.9324748333};
test_output[2956] = '{137.759899455};
############ END DEBUG ############*/
test_input[23656:23663] = '{32'hc112990b, 32'hc18fb26a, 32'h41b3d332, 32'hc2b960f8, 32'h42a69f48, 32'h411e875b, 32'h42828ea6, 32'hc280f97f};
test_label[2957] = '{32'h42a69f48};
test_output[2957] = '{32'h327d48f3};
/*############ DEBUG ############
test_input[23656:23663] = '{-9.16236417622, -17.9621170213, 22.4781232977, -92.689394236, 83.3110967123, 9.90804531064, 65.2786077346, -64.4872998757};
test_label[2957] = '{83.3110967123};
test_output[2957] = '{1.47431247187e-08};
############ END DEBUG ############*/
test_input[23664:23671] = '{32'hc1209175, 32'h41c04631, 32'h41a36f98, 32'h4222fab1, 32'hc2bcf8ac, 32'hc1c7f63e, 32'h424c07ff, 32'h42c2c3dc};
test_label[2958] = '{32'h42c2c3dc};
test_output[2958] = '{32'h80000000};
/*############ DEBUG ############
test_input[23664:23671] = '{-10.0355118855, 24.0342729972, 20.4294898085, 40.7448139637, -94.4856860122, -24.9952351761, 51.007807459, 97.3825348703};
test_label[2958] = '{97.3825348703};
test_output[2958] = '{-0.0};
############ END DEBUG ############*/
test_input[23672:23679] = '{32'h4182b137, 32'hc203ab9d, 32'h42b8220b, 32'hc288ebf8, 32'h424e4e0c, 32'h42abf1ba, 32'hc2a8ecc8, 32'hc2705041};
test_label[2959] = '{32'h42b8220b};
test_output[2959] = '{32'h3b13a6de};
/*############ DEBUG ############
test_input[23672:23679] = '{16.3365302498, -32.91759016, 92.0664904994, -68.4608777408, 51.5762195384, 85.9721192414, -84.4624662367, -60.078371708};
test_label[2959] = '{92.0664904994};
test_output[2959] = '{0.00225298795567};
############ END DEBUG ############*/
test_input[23680:23687] = '{32'h421b3204, 32'h42405f60, 32'hc2a4e4e6, 32'hc2575008, 32'hc261ccc8, 32'hc1db2766, 32'hc2a4f10a, 32'hc2a5941c};
test_label[2960] = '{32'hc1db2766};
test_output[2960] = '{32'h4296f995};
/*############ DEBUG ############
test_input[23680:23687] = '{38.7988438904, 48.0931387758, -82.447064585, -53.8281544947, -56.4499813446, -27.3942366135, -82.4707788239, -82.7892742138};
test_label[2960] = '{-27.3942366135};
test_output[2960] = '{75.4874673324};
############ END DEBUG ############*/
test_input[23688:23695] = '{32'hc277d797, 32'hc21059c0, 32'h429933ae, 32'hc2b2c3c7, 32'h428c00fa, 32'hc2873e70, 32'hbf023fea, 32'h41e4343f};
test_label[2961] = '{32'hc21059c0};
test_output[2961] = '{32'h42e16140};
/*############ DEBUG ############
test_input[23688:23695] = '{-61.9605378106, -36.0876455675, 76.6009348954, -89.3823769994, 70.0019070767, -67.6219489659, -0.508787771514, 28.5255112987};
test_label[2961] = '{-36.0876455675};
test_output[2961] = '{112.689941228};
############ END DEBUG ############*/
test_input[23696:23703] = '{32'h428109f4, 32'hc2c5067b, 32'hc2b60db6, 32'h41d9322c, 32'hbf26752b, 32'hc2af10da, 32'hc29e5139, 32'h41b7d56a};
test_label[2962] = '{32'hc2b60db6};
test_output[2962] = '{32'h431b8bd5};
/*############ DEBUG ############
test_input[23696:23703] = '{64.5194432005, -98.5126606144, -91.0267820421, 27.1494972974, -0.650225354867, -87.532916609, -79.1586342826, 22.9792051367};
test_label[2962] = '{-91.0267820421};
test_output[2962] = '{155.546225243};
############ END DEBUG ############*/
test_input[23704:23711] = '{32'hc29cecb3, 32'h40d13385, 32'hc126f8e4, 32'h42b4558b, 32'hc2bde20b, 32'hc291eacd, 32'hc2b621fb, 32'h42bc38c2};
test_label[2963] = '{32'hc29cecb3};
test_output[2963] = '{32'h432c97a4};
/*############ DEBUG ############
test_input[23704:23711] = '{-78.4623052574, 6.53753887444, -10.4357642339, 90.1670785183, -94.9414883694, -72.9585987333, -91.0663669479, 94.1108514989};
test_label[2963] = '{-78.4623052574};
test_output[2963] = '{172.592346426};
############ END DEBUG ############*/
test_input[23712:23719] = '{32'h4294464a, 32'h424ac863, 32'hc205d41d, 32'hc2047b44, 32'h428cef96, 32'hc286c704, 32'h428bcc1e, 32'hc2a68f9d};
test_label[2964] = '{32'hc205d41d};
test_output[2964] = '{32'h42d74463};
/*############ DEBUG ############
test_input[23712:23719] = '{74.1372842556, 50.6956904434, -33.4571413428, -33.1203780806, 70.4679442423, -67.3887034524, 69.8986677533, -83.2804931721};
test_label[2964] = '{-33.4571413428};
test_output[2964] = '{107.633570182};
############ END DEBUG ############*/
test_input[23720:23727] = '{32'h429c9258, 32'hc196244d, 32'hc148c1b1, 32'hc2a2a280, 32'h4285ddf2, 32'h425a0f03, 32'hbf8c96f0, 32'hc28712f4};
test_label[2965] = '{32'hc2a2a280};
test_output[2965] = '{32'h431f9a6d};
/*############ DEBUG ############
test_input[23720:23727] = '{78.2858306517, -18.7677245061, -12.5472881348, -81.3173799565, 66.9334881795, 54.5146583784, -1.09835624619, -67.5370178202};
test_label[2965] = '{-81.3173799565};
test_output[2965] = '{159.60322235};
############ END DEBUG ############*/
test_input[23728:23735] = '{32'h422d5f8a, 32'hc2815357, 32'hc0fe11e2, 32'hc1ec1d9f, 32'hc1e7296d, 32'h4298d1f9, 32'h4150f844, 32'hc2a23522};
test_label[2966] = '{32'h4298d1f9};
test_output[2966] = '{32'h279c0000};
/*############ DEBUG ############
test_input[23728:23735] = '{43.3433010679, -64.6627693914, -7.9396829581, -29.5144628178, -28.8952281572, 76.4101002753, 13.0606121367, -81.1037719994};
test_label[2966] = '{76.4101002753};
test_output[2966] = '{4.32986979604e-15};
############ END DEBUG ############*/
test_input[23736:23743] = '{32'h413abbde, 32'hc2ac03a0, 32'hc1e703e9, 32'hc2ad5c51, 32'hc22faccb, 32'h4162fb8b, 32'h42c39d5a, 32'hc22cbca1};
test_label[2967] = '{32'h413abbde};
test_output[2967] = '{32'h42ac45de};
/*############ DEBUG ############
test_input[23736:23743] = '{11.6708655444, -86.0070820444, -28.8769096633, -86.6803069414, -43.9187445956, 14.1864115202, 97.8073256098, -43.1842060089};
test_label[2967] = '{11.6708655444};
test_output[2967] = '{86.1364600653};
############ END DEBUG ############*/
test_input[23744:23751] = '{32'h42763458, 32'h3f36d474, 32'h424df150, 32'hc1753851, 32'h429de85a, 32'hc1e21099, 32'hc108c959, 32'h41bdac5b};
test_label[2968] = '{32'hc1e21099};
test_output[2968] = '{32'h42d66c81};
/*############ DEBUG ############
test_input[23744:23751] = '{61.5511183245, 0.714179302128, 51.4856550478, -15.3262489595, 78.9538143185, -28.2581039249, -8.54915679421, 23.7091571632};
test_label[2968] = '{-28.2581039249};
test_output[2968] = '{107.211918271};
############ END DEBUG ############*/
test_input[23752:23759] = '{32'hc2a65a04, 32'hc2214509, 32'hc0943ece, 32'h4250000b, 32'hc23ba2d8, 32'h4298797a, 32'h3fb28d6f, 32'h40a05e0b};
test_label[2969] = '{32'hc2a65a04};
test_output[2969] = '{32'h431f69bf};
/*############ DEBUG ############
test_input[23752:23759] = '{-83.1758137726, -40.3174155382, -4.63266674772, 52.000040119, -46.9090281981, 76.2372573114, 1.39494121304, 5.01147989554};
test_label[2969] = '{-83.1758137726};
test_output[2969] = '{159.413071084};
############ END DEBUG ############*/
test_input[23760:23767] = '{32'hc23700a1, 32'h4154c086, 32'h40625641, 32'h42b05823, 32'h42bb7756, 32'hc1cb1a2e, 32'hc2c79eb3, 32'hc21434f9};
test_label[2970] = '{32'hc23700a1};
test_output[2970] = '{32'h430b7ccf};
/*############ DEBUG ############
test_input[23760:23767] = '{-45.7506138512, 13.29700264, 3.5365146361, 88.1721437413, 93.7330753845, -25.3877832092, -99.8099621815, -37.0517314169};
test_label[2970] = '{-45.7506138512};
test_output[2970] = '{139.487527054};
############ END DEBUG ############*/
test_input[23768:23775] = '{32'hc299e8cb, 32'h42a609fe, 32'hc23008e1, 32'hc2727606, 32'hc23b9a68, 32'hc2aa3d28, 32'hc2a778d4, 32'hc0a948af};
test_label[2971] = '{32'hc23008e1};
test_output[2971] = '{32'h42fe0e6e};
/*############ DEBUG ############
test_input[23768:23775] = '{-76.9546754238, 83.0195127044, -44.0086696288, -60.6152582486, -46.9007877067, -85.1194483682, -83.7359943428, -5.29012258552};
test_label[2971] = '{-44.0086696288};
test_output[2971] = '{127.028182333};
############ END DEBUG ############*/
test_input[23776:23783] = '{32'h417ca494, 32'h4106de02, 32'h42915479, 32'hc2104c59, 32'hc2a9362e, 32'h4227b821, 32'hc262fff6, 32'h4207a99d};
test_label[2972] = '{32'hc262fff6};
test_output[2972] = '{32'h43016a3a};
/*############ DEBUG ############
test_input[23776:23783] = '{15.7901804597, 8.42920157286, 72.6649882939, -36.0745585334, -84.6058205223, 41.9298149568, -56.749963628, 33.915638319};
test_label[2972] = '{-56.749963628};
test_output[2972] = '{129.414951922};
############ END DEBUG ############*/
test_input[23784:23791] = '{32'h4219409e, 32'h3fd18504, 32'hc1fcc63e, 32'h42899e42, 32'h422b7211, 32'h422af581, 32'hc25a8e49, 32'hc28ed123};
test_label[2973] = '{32'h42899e42};
test_output[2973] = '{32'h2d339180};
/*############ DEBUG ############
test_input[23784:23791] = '{38.3131014948, 1.63687181893, -31.59679702, 68.8090952566, 42.8613923382, 42.7397488706, -54.6389507318, -71.4084689989};
test_label[2973] = '{68.8090952566};
test_output[2973] = '{1.02072794662e-11};
############ END DEBUG ############*/
test_input[23792:23799] = '{32'hc26f2116, 32'hc25235ef, 32'hc1c8d23d, 32'hc16120ba, 32'h41e848f1, 32'hc2674838, 32'h4140cc34, 32'h42c0dfb5};
test_label[2974] = '{32'h41e848f1};
test_output[2974] = '{32'h4286cd79};
/*############ DEBUG ############
test_input[23792:23799] = '{-59.7823102636, -52.5526683183, -25.1026559158, -14.0704901137, 29.0356152705, -57.8205278859, 12.0498541248, 96.4369312464};
test_label[2974] = '{29.0356152705};
test_output[2974] = '{67.4013159759};
############ END DEBUG ############*/
test_input[23800:23807] = '{32'h40c8a875, 32'h425af9cb, 32'hc1cb65fb, 32'hc297ebfd, 32'h41d59eb8, 32'h4104516f, 32'hc21fd70e, 32'h424770e3};
test_label[2975] = '{32'h4104516f};
test_output[2975] = '{32'h4239ed28};
/*############ DEBUG ############
test_input[23800:23807] = '{6.27056340597, 54.7439379787, -25.4247960892, -75.9609168841, 26.7024987978, 8.26988127055, -39.9600148157, 49.8602409744};
test_label[2975] = '{8.26988127055};
test_output[2975] = '{46.4815971868};
############ END DEBUG ############*/
test_input[23808:23815] = '{32'hc1096a15, 32'hc11f97db, 32'h41c23c63, 32'h424914d0, 32'h4264ee89, 32'h423a4277, 32'hc2be4c46, 32'h42bbf528};
test_label[2976] = '{32'hc2be4c46};
test_output[2976] = '{32'h433d20b7};
/*############ DEBUG ############
test_input[23808:23815] = '{-8.58839876091, -9.97457440683, 24.2794848355, 50.270323737, 57.2329461658, 46.5649053658, -95.1489685125, 93.9788173505};
test_label[2976] = '{-95.1489685125};
test_output[2976] = '{189.127785863};
############ END DEBUG ############*/
test_input[23816:23823] = '{32'hc1d1556c, 32'h428a7e07, 32'hc1da1edc, 32'hc2904f5d, 32'hc294f3a6, 32'hc2a66e99, 32'h4218b741, 32'hc2a45414};
test_label[2977] = '{32'h4218b741};
test_output[2977] = '{32'h41f8899a};
/*############ DEBUG ############
test_input[23816:23823] = '{-26.166709952, 69.2461468985, -27.2650685418, -72.1550045591, -74.4758721586, -83.2160096872, 38.1789590644, -82.1642131003};
test_label[2977] = '{38.1789590644};
test_output[2977] = '{31.0671878341};
############ END DEBUG ############*/
test_input[23824:23831] = '{32'hc22974b4, 32'hc21ac032, 32'h40543b71, 32'hc2a7dc97, 32'h420b4542, 32'hc0a73a7b, 32'hc2a34b96, 32'h4242fd4b};
test_label[2978] = '{32'h420b4542};
test_output[2978] = '{32'h415ee027};
/*############ DEBUG ############
test_input[23824:23831] = '{-42.3639663569, -38.6876906815, 3.31612807172, -83.9308359083, 34.8176335681, -5.22588891447, -81.6476265786, 48.7473577988};
test_label[2978] = '{34.8176335681};
test_output[2978] = '{13.9297251228};
############ END DEBUG ############*/
test_input[23832:23839] = '{32'hc2221a1a, 32'hc24d8a39, 32'hc285fb78, 32'h41814313, 32'hc1e18739, 32'h4226dc2f, 32'h40e87274, 32'h41c60a68};
test_label[2979] = '{32'hc24d8a39};
test_output[2979] = '{32'h42ba3334};
/*############ DEBUG ############
test_input[23832:23839] = '{-40.5254881882, -51.3849834965, -66.9911481629, 16.1577505234, -28.1910272837, 41.7150212457, 7.26397143134, 24.7550803679};
test_label[2979] = '{-51.3849834965};
test_output[2979] = '{93.1000047853};
############ END DEBUG ############*/
test_input[23840:23847] = '{32'hc1ea751c, 32'hc1fd8a8f, 32'hc18a0fe5, 32'h4241b84f, 32'hc208de72, 32'hc2a42eb7, 32'hc1e9850e, 32'hc2aa7c8f};
test_label[2980] = '{32'hc1ea751c};
test_output[2980] = '{32'h429b796e};
/*############ DEBUG ############
test_input[23840:23847] = '{-29.3071819934, -31.6926549733, -17.2577613586, 48.4299883199, -34.2172335661, -82.0912403194, -29.1899688003, -85.243276317};
test_label[2980] = '{-29.3071819934};
test_output[2980] = '{77.7371703133};
############ END DEBUG ############*/
test_input[23848:23855] = '{32'hc1a0ed05, 32'h420903b9, 32'h42493ecb, 32'hc19f0f57, 32'h41980f33, 32'h42bea509, 32'h42ac4037, 32'h425ca0be};
test_label[2981] = '{32'h41980f33};
test_output[2981] = '{32'h4298a149};
/*############ DEBUG ############
test_input[23848:23855] = '{-20.1157327634, 34.2536371879, 50.3113205032, -19.8824901061, 19.0074215086, 95.3223334659, 86.1254214007, 55.1569739364};
test_label[2981] = '{19.0074215086};
test_output[2981] = '{76.3150133041};
############ END DEBUG ############*/
test_input[23856:23863] = '{32'hc26b245a, 32'h42b04343, 32'h422fe2c2, 32'h42bfdf8a, 32'h42b1f43b, 32'hc212f7c4, 32'h42a70ea7, 32'hc1aebaf9};
test_label[2982] = '{32'h422fe2c2};
test_output[2982] = '{32'h424fddb7};
/*############ DEBUG ############
test_input[23856:23863] = '{-58.7855001013, 88.1313711116, 43.9714444624, 95.9366011469, 88.9770139403, -36.7419572467, 83.5286153045, -21.8412961765};
test_label[2982] = '{43.9714444624};
test_output[2982] = '{51.9665169308};
############ END DEBUG ############*/
test_input[23864:23871] = '{32'h4297ac1f, 32'hc21311c1, 32'hc2643e65, 32'h428b66e7, 32'hc20a1e39, 32'hc299e631, 32'hbf859e87, 32'h42b6c3f2};
test_label[2983] = '{32'hc21311c1};
test_output[2983] = '{32'h43002669};
/*############ DEBUG ############
test_input[23864:23871] = '{75.8361745302, -36.7673386655, -57.0609323143, 69.7009810712, -34.5295124762, -76.9495942035, -1.04390040721, 91.3827049059};
test_label[2983] = '{-36.7673386655};
test_output[2983] = '{128.150043749};
############ END DEBUG ############*/
test_input[23872:23879] = '{32'hc2b81dda, 32'h4279f075, 32'hc27ed389, 32'h41073196, 32'hc2b8f67f, 32'hc2210ab7, 32'hc2c5b28d, 32'h4173001d};
test_label[2984] = '{32'h41073196};
test_output[2984] = '{32'h4258240f};
/*############ DEBUG ############
test_input[23872:23879] = '{-92.0583023076, 62.4848210043, -63.7065763969, 8.44960593489, -92.4814380213, -40.2604644519, -98.8487303737, 15.1875279115};
test_label[2984] = '{8.44960593489};
test_output[2984] = '{54.0352150694};
############ END DEBUG ############*/
test_input[23880:23887] = '{32'hc055d1d3, 32'h428304ad, 32'hc1916683, 32'h425d4dcc, 32'h413d2285, 32'h428e72ae, 32'h4261193a, 32'h4297e746};
test_label[2985] = '{32'h4261193a};
test_output[2985] = '{32'h419d7cba};
/*############ DEBUG ############
test_input[23880:23887] = '{-3.34093159384, 65.5091332799, -18.1750544422, 55.3259716923, 11.8209274236, 71.2239843048, 56.274636502, 75.9517021288};
test_label[2985] = '{56.274636502};
test_output[2985] = '{19.6859022741};
############ END DEBUG ############*/
test_input[23888:23895] = '{32'h429532f1, 32'h41f924b7, 32'h4245619b, 32'hc1a92f20, 32'h42bdf968, 32'h42afd992, 32'h42c12663, 32'h425a4539};
test_label[2986] = '{32'h425a4539};
test_output[2986] = '{32'h4228c61d};
/*############ DEBUG ############
test_input[23888:23895] = '{74.5994949197, 31.1429263161, 49.3453175526, -21.1480097063, 94.9871236318, 87.9249445467, 96.5749739875, 54.5676020196};
test_label[2986] = '{54.5676020196};
test_output[2986] = '{42.1934693646};
############ END DEBUG ############*/
test_input[23896:23903] = '{32'h40a55dc1, 32'hc1aef9bb, 32'hc23baf3b, 32'h429c971d, 32'h41e544b3, 32'hc20f60cc, 32'h4170b1d8, 32'h42a95418};
test_label[2987] = '{32'h4170b1d8};
test_output[2987] = '{32'h428b3ebe};
/*############ DEBUG ############
test_input[23896:23903] = '{5.16769473914, -21.8719386269, -46.9211236501, 78.2951421953, 28.6585440195, -35.8445275297, 15.0434188187, 84.664247219};
test_label[2987] = '{15.0434188187};
test_output[2987] = '{69.6225406258};
############ END DEBUG ############*/
test_input[23904:23911] = '{32'hc2ba01fd, 32'hc0be071e, 32'h4116aa53, 32'h408d955f, 32'hc265aba3, 32'h42a75037, 32'h42a3d6f7, 32'hc2a19132};
test_label[2988] = '{32'h42a75037};
test_output[2988] = '{32'h3e26143d};
/*############ DEBUG ############
test_input[23904:23911] = '{-93.003886197, -5.93836876122, 9.41658288738, 4.42448355308, -57.4176128289, 83.6566722806, 81.9198534235, -80.7835824885};
test_label[2988] = '{83.6566722806};
test_output[2988] = '{0.162186572637};
############ END DEBUG ############*/
test_input[23912:23919] = '{32'h422306e7, 32'h4273dfa8, 32'hc1bb64e8, 32'h41beeeea, 32'h41ea85a4, 32'hc2bb8a97, 32'h42c4a313, 32'h42820855};
test_label[2989] = '{32'hc2bb8a97};
test_output[2989] = '{32'h434016d5};
/*############ DEBUG ############
test_input[23912:23919] = '{40.7567423175, 60.9684159292, -23.4242700733, 23.8666575263, 29.3152542846, -93.7706820558, 98.3185022109, 65.0162733141};
test_label[2989] = '{-93.7706820558};
test_output[2989] = '{192.089184267};
############ END DEBUG ############*/
test_input[23920:23927] = '{32'hc2b23639, 32'hc1566149, 32'h42a063c0, 32'hc20868cb, 32'h42164540, 32'h416751ad, 32'h413a19ce, 32'hc1524699};
test_label[2990] = '{32'hc1566149};
test_output[2990] = '{32'h42bb2fe9};
/*############ DEBUG ############
test_input[23920:23927] = '{-89.1059027392, -13.3987517246, 80.1948248035, -34.1023376887, 37.5676274289, 14.4574401942, 11.6312995844, -13.1422354786};
test_label[2990] = '{-13.3987517246};
test_output[2990] = '{93.5935765281};
############ END DEBUG ############*/
test_input[23928:23935] = '{32'h42558256, 32'h41d6be85, 32'h4185d3be, 32'hc180a453, 32'h42c40158, 32'hc2c52a8f, 32'h41da5546, 32'h425cce4d};
test_label[2991] = '{32'h42558256};
test_output[2991] = '{32'h4232805b};
/*############ DEBUG ############
test_input[23928:23935] = '{53.3772796286, 26.8430263386, 16.7283895432, -16.0802373685, 98.0026273852, -98.583124243, 27.2916366395, 55.2014640604};
test_label[2991] = '{53.3772796286};
test_output[2991] = '{44.6253477566};
############ END DEBUG ############*/
test_input[23936:23943] = '{32'hc2a4f2d5, 32'h4104192e, 32'h41ce5084, 32'hc24f60c8, 32'hc2366ca1, 32'hc23e7f5d, 32'h41af6f55, 32'hc21a841d};
test_label[2992] = '{32'hc21a841d};
test_output[2992] = '{32'h4280e0dc};
/*############ DEBUG ############
test_input[23936:23943] = '{-82.4742849012, 8.25614782251, 25.7893134181, -51.844511225, -45.6060841787, -47.6243768408, 21.9293618797, -38.6290178777};
test_label[2992] = '{-38.6290178777};
test_output[2992] = '{64.4391814574};
############ END DEBUG ############*/
test_input[23944:23951] = '{32'hc2adf438, 32'hc127e30f, 32'hc154c453, 32'hc253e061, 32'hc003ae07, 32'hc2bfe729, 32'hc21fb124, 32'hc2281aea};
test_label[2993] = '{32'hc003ae07};
test_output[2993] = '{32'h397152d0};
/*############ DEBUG ############
test_input[23944:23951] = '{-86.9769897882, -10.4929341235, -13.2979305865, -52.9691182201, -2.05749682274, -95.9514859806, -39.9229895025, -42.0262839075};
test_label[2993] = '{-2.05749682274};
test_output[2993] = '{0.000230144014899};
############ END DEBUG ############*/
test_input[23952:23959] = '{32'h42b824ea, 32'hc1930c87, 32'h42984916, 32'hc2153387, 32'h4229aba0, 32'hc231b5d9, 32'hc2a1b38a, 32'hc18753d5};
test_label[2994] = '{32'hc2153387};
test_output[2994] = '{32'h43015f57};
/*############ DEBUG ############
test_input[23952:23959] = '{92.0720966086, -18.3811166912, 76.1427434332, -37.3003189316, 42.4176017853, -44.4275855817, -80.85066042, -16.9159335586};
test_label[2994] = '{-37.3003189316};
test_output[2994] = '{129.372415661};
############ END DEBUG ############*/
test_input[23960:23967] = '{32'h4280c1dd, 32'h42735073, 32'h4299cacf, 32'hc1493fcb, 32'hc28842b4, 32'hc2be4523, 32'hc2c50843, 32'hc1c2f0df};
test_label[2995] = '{32'hc28842b4};
test_output[2995] = '{32'h431106c2};
/*############ DEBUG ############
test_input[23960:23967] = '{64.3786396262, 60.8285639653, 76.8961083573, -12.5780742774, -68.1302818297, -95.1350345418, -98.5161342816, -24.3676126323};
test_label[2995] = '{-68.1302818297};
test_output[2995] = '{145.026393954};
############ END DEBUG ############*/
test_input[23968:23975] = '{32'hc25dbe11, 32'hc1d2975c, 32'hc1a4153f, 32'hc288db77, 32'hc26b182d, 32'h4209b43d, 32'hc0923ac5, 32'hc1f4ef63};
test_label[2996] = '{32'hc1f4ef63};
test_output[2996] = '{32'h428215f8};
/*############ DEBUG ############
test_input[23968:23975] = '{-55.4356119184, -26.3239067336, -20.5103742116, -68.4286423175, -58.7736087549, 34.4260155423, -4.569673903, -30.6168888703};
test_label[2996] = '{-30.6168888703};
test_output[2996] = '{65.0429044126};
############ END DEBUG ############*/
test_input[23976:23983] = '{32'h42964563, 32'h40973ab0, 32'hc24d97c8, 32'h40f1c030, 32'hc25988fd, 32'hc296a319, 32'h42be7346, 32'h4165cf3e};
test_label[2997] = '{32'h40f1c030};
test_output[2997] = '{32'h42af5743};
/*############ DEBUG ############
test_input[23976:23983] = '{75.1355239672, 4.72591415669, -51.3982225285, 7.55471034534, -54.3837765462, -75.3185523014, 95.2251463437, 14.3630964621};
test_label[2997] = '{7.55471034534};
test_output[2997] = '{87.6704360002};
############ END DEBUG ############*/
test_input[23984:23991] = '{32'h4286b0f6, 32'h41de1cd5, 32'h42b3c25a, 32'h425184a0, 32'hc22ec56f, 32'h41467015, 32'hc01115ba, 32'h42805242};
test_label[2998] = '{32'h4286b0f6};
test_output[2998] = '{32'h41b44593};
/*############ DEBUG ############
test_input[23984:23991] = '{67.3456236473, 27.7640780535, 89.8795949047, 52.3795182345, -43.6928064344, 12.4023641848, -2.26695098876, 64.1606632487};
test_label[2998] = '{67.3456236473};
test_output[2998] = '{22.5339712576};
############ END DEBUG ############*/
test_input[23992:23999] = '{32'hc2a9c660, 32'h423d622b, 32'h3f8f788e, 32'hc28b5d2b, 32'hc1dd8297, 32'h4198d098, 32'h423e4dc7, 32'h427aba02};
test_label[2999] = '{32'hc28b5d2b};
test_output[2999] = '{32'h43045d16};
/*############ DEBUG ############
test_input[23992:23999] = '{-84.8874498715, 47.3458666472, 1.12086658799, -69.6819702518, -27.6887651411, 19.1018515978, 47.5759529637, 62.6816470358};
test_label[2999] = '{-69.6819702518};
test_output[2999] = '{132.363617781};
############ END DEBUG ############*/
test_input[24000:24007] = '{32'hc26fdf00, 32'hc007dabf, 32'h428885a1, 32'hc2b962b7, 32'hc2bba09b, 32'hc244d721, 32'h41fda2a9, 32'h42c7cd9d};
test_label[3000] = '{32'hc244d721};
test_output[3000] = '{32'h43151c97};
/*############ DEBUG ############
test_input[24000:24007] = '{-59.9677731812, -2.1227262113, 68.260990578, -92.6928000444, -93.8136832172, -49.2100855321, 31.7044246236, 99.901587441};
test_label[3000] = '{-49.2100855321};
test_output[3000] = '{149.111672973};
############ END DEBUG ############*/
test_input[24008:24015] = '{32'h4205e977, 32'hc1ac94e6, 32'hc1e451ef, 32'hc10be750, 32'h42392c1d, 32'h4104863d, 32'h41837d4e, 32'hc228d99a};
test_label[3001] = '{32'h41837d4e};
test_output[3001] = '{32'h41eedaee};
/*############ DEBUG ############
test_input[24008:24015] = '{33.477993125, -21.572704525, -28.540007401, -8.74397265496, 46.2930799637, 8.28277328421, 16.4361837197, -42.2125031015};
test_label[3001] = '{16.4361837197};
test_output[3001] = '{29.8568989634};
############ END DEBUG ############*/
test_input[24016:24023] = '{32'hc191981b, 32'hc1bae645, 32'h428c49ab, 32'h41d3b1a3, 32'h425fa3d7, 32'h410cd7ea, 32'hc28be1b4, 32'h424b86b8};
test_label[3002] = '{32'h425fa3d7};
test_output[3002] = '{32'h4163be00};
/*############ DEBUG ############
test_input[24016:24023] = '{-18.199269725, -23.3624364486, 70.1438845386, 26.4617375933, 55.9099980939, 8.80271339158, -69.9408297617, 50.8815602428};
test_label[3002] = '{55.9099980939};
test_output[3002] = '{14.2338871071};
############ END DEBUG ############*/
test_input[24024:24031] = '{32'h41a1371d, 32'hc2af0b51, 32'h42bb7546, 32'h42b5db71, 32'h4220b646, 32'hc19115d1, 32'h41bfd437, 32'h428a5b6a};
test_label[3003] = '{32'h41bfd437};
test_output[3003] = '{32'h428b9e6f};
/*############ DEBUG ############
test_input[24024:24031] = '{20.1519104989, -87.522101822, 93.7290525428, 90.9285950594, 40.1780031125, -18.1356523837, 23.9786205249, 69.1785397652};
test_label[3003] = '{23.9786205249};
test_output[3003] = '{69.8094386251};
############ END DEBUG ############*/
test_input[24032:24039] = '{32'hc23ca43d, 32'hc18578ee, 32'hc27035d5, 32'hc248f896, 32'hc198990f, 32'h419214f0, 32'hc28a6a40, 32'hc178df66};
test_label[3004] = '{32'hc27035d5};
test_output[3004] = '{32'h429ca027};
/*############ DEBUG ############
test_input[24032:24039] = '{-47.160388981, -16.6840470091, -60.0525719905, -50.2427612809, -19.074736323, 18.2602230565, -69.2075162275, -15.5545402794};
test_label[3004] = '{-60.0525719905};
test_output[3004] = '{78.312795047};
############ END DEBUG ############*/
test_input[24040:24047] = '{32'h4256e59f, 32'h40b56dba, 32'h42bc4558, 32'hc2119851, 32'h41de2f6d, 32'hc22818ed, 32'hc225fa31, 32'h42831279};
test_label[3005] = '{32'h41de2f6d};
test_output[3005] = '{32'h4284b97c};
/*############ DEBUG ############
test_input[24040:24047] = '{53.7242385786, 5.66964442663, 94.1354334586, -36.3987450268, 27.7731571149, -42.0243424897, -41.4943285449, 65.5360825405};
test_label[3005] = '{27.7731571149};
test_output[3005] = '{66.3622763437};
############ END DEBUG ############*/
test_input[24048:24055] = '{32'h4282243b, 32'h42a75416, 32'h427ea361, 32'hc2c602c4, 32'hc259d6b8, 32'h42b3b526, 32'hc2bb6136, 32'hc1580e8e};
test_label[3006] = '{32'h427ea361};
test_output[3006] = '{32'h41d19207};
/*############ DEBUG ############
test_input[24048:24055] = '{65.0707630496, 83.6642265658, 63.6595481778, -99.0054000571, -54.4596862681, 89.8538020786, -93.6898681201, -13.5035534286};
test_label[3006] = '{63.6595481778};
test_output[3006] = '{26.196302498};
############ END DEBUG ############*/
test_input[24056:24063] = '{32'hc2a22fa4, 32'hc126cd40, 32'hc2b9752e, 32'h420645f4, 32'hc2b66718, 32'hc2b33840, 32'hc192f63a, 32'h4108ef4b};
test_label[3007] = '{32'h4108ef4b};
test_output[3007] = '{32'h41c81442};
/*############ DEBUG ############
test_input[24056:24063] = '{-81.0930511293, -10.4251102808, -92.728863433, 33.5683119442, -91.2013555539, -89.6098662655, -18.3702283311, 8.5584211869};
test_label[3007] = '{8.5584211869};
test_output[3007] = '{25.0098907573};
############ END DEBUG ############*/
test_input[24064:24071] = '{32'h415cf0fb, 32'hc2b882e1, 32'h4209bb55, 32'h4251ca52, 32'h4267d5d9, 32'h4134c326, 32'h429b8c62, 32'hc2898a47};
test_label[3008] = '{32'h4267d5d9};
test_output[3008] = '{32'h419e85d5};
/*############ DEBUG ############
test_input[24064:24071] = '{13.8088328194, -92.2556218158, 34.4329398479, 52.4475775579, 57.9588372908, 11.2976441206, 77.7741847516, -68.7700723365};
test_label[3008] = '{57.9588372908};
test_output[3008] = '{19.8153474633};
############ END DEBUG ############*/
test_input[24072:24079] = '{32'h427a2549, 32'h42c0f470, 32'h42bc68d8, 32'h40aa5e16, 32'h42a5274f, 32'hc18e0437, 32'hc223c9c3, 32'hc21ad10f};
test_label[3009] = '{32'h42a5274f};
test_output[3009] = '{32'h415ffab6};
/*############ DEBUG ############
test_input[24072:24079] = '{62.5364121138, 96.4774139861, 94.204769723, 5.32398523226, 82.576775979, -17.7520571629, -40.9470315048, -38.704160569};
test_label[3009] = '{82.576775979};
test_output[3009] = '{13.9987082606};
############ END DEBUG ############*/
test_input[24080:24087] = '{32'hc2aebbf8, 32'hc2994625, 32'h41657b0d, 32'hc293127e, 32'hc2bb273e, 32'hc2923e2e, 32'h420a2258, 32'hc2ae1afe};
test_label[3010] = '{32'hc2994625};
test_output[3010] = '{32'h42de5751};
/*############ DEBUG ############
test_input[24080:24087] = '{-87.3671287958, -76.6369994936, 14.3425416165, -73.536116057, -93.5766415547, -73.1214413372, 34.5335399913, -87.0527220994};
test_label[3010] = '{-76.6369994936};
test_output[3010] = '{111.170539487};
############ END DEBUG ############*/
test_input[24088:24095] = '{32'h4225f70b, 32'hc29c70a7, 32'h4242f328, 32'h4220da2c, 32'hc25e8ae4, 32'h42471a63, 32'hc1c50f8f, 32'h42534de2};
test_label[3011] = '{32'h4242f328};
test_output[3011] = '{32'h4084d2f1};
/*############ DEBUG ############
test_input[24088:24095] = '{41.4912532378, -78.2200208254, 48.7374590589, 40.2130565822, -55.6356336605, 49.7757688595, -24.6325972212, 52.826057488};
test_label[3011] = '{48.7374590589};
test_output[3011] = '{4.15074964658};
############ END DEBUG ############*/
test_input[24096:24103] = '{32'h42a19faf, 32'h4289227f, 32'h41076a47, 32'hc0742aac, 32'h42702641, 32'hc18cfe38, 32'h412e6d73, 32'hc015ce13};
test_label[3012] = '{32'h42a19faf};
test_output[3012] = '{32'h36a17a52};
/*############ DEBUG ############
test_input[24096:24103] = '{80.8118843355, 68.5673775122, 8.46344662089, -3.81510438025, 60.037357499, -17.6241301901, 10.9017211649, -2.34070269706};
test_label[3012] = '{80.8118843355};
test_output[3012] = '{4.81241366592e-06};
############ END DEBUG ############*/
test_input[24104:24111] = '{32'hc2adfa11, 32'hc14ca653, 32'hc23f813e, 32'hc2bfec6b, 32'hc2a76023, 32'hc27d9272, 32'hc29d4e26, 32'h40ded25d};
test_label[3013] = '{32'hc27d9272};
test_output[3013] = '{32'h428cb65f};
/*############ DEBUG ############
test_input[24104:24111] = '{-86.9884086915, -12.7906065146, -47.8762116888, -95.9617540691, -83.6877708164, -63.3930123076, -78.6526329803, 6.96317894457};
test_label[3013] = '{-63.3930123076};
test_output[3013] = '{70.3561912548};
############ END DEBUG ############*/
test_input[24112:24119] = '{32'h42046573, 32'h42b05d4e, 32'h42b22ec8, 32'h4282033a, 32'h42ab785f, 32'h428ef5a9, 32'hc205bdc2, 32'hc28c306e};
test_label[3014] = '{32'h42b05d4e};
test_output[3014] = '{32'h3fa2d79b};
/*############ DEBUG ############
test_input[24112:24119] = '{33.0990721726, 88.1822343964, 89.0913679334, 65.0063053916, 85.7351006074, 71.4798035736, -33.4353097271, -70.094592237};
test_label[3014] = '{88.1822343964};
test_output[3014] = '{1.27220480944};
############ END DEBUG ############*/
test_input[24120:24127] = '{32'hc257bfba, 32'h411c8615, 32'h42beece2, 32'h41ffdc8f, 32'h42647495, 32'h4231f364, 32'h42779e44, 32'hc22bfd88};
test_label[3015] = '{32'h42779e44};
test_output[3015] = '{32'h42063b80};
/*############ DEBUG ############
test_input[24120:24127] = '{-53.9372331708, 9.78273519193, 95.4626646075, 31.9826948798, 57.1138491504, 44.4876855153, 61.9045573791, -42.9975901365};
test_label[3015] = '{61.9045573791};
test_output[3015] = '{33.5581072284};
############ END DEBUG ############*/
test_input[24128:24135] = '{32'h4293dfb4, 32'h42591d70, 32'h42c5a5e8, 32'h41e0679d, 32'hc281f279, 32'h42af5b75, 32'h428e967e, 32'hc1466a1b};
test_label[3016] = '{32'h42af5b75};
test_output[3016] = '{32'h413253ad};
/*############ DEBUG ############
test_input[24128:24135] = '{73.9369223532, 54.2787489415, 98.8240379556, 28.0505921876, -64.9735770656, 87.6786234118, 71.2939337213, -12.4009042647};
test_label[3016] = '{87.6786234118};
test_output[3016] = '{11.1454289851};
############ END DEBUG ############*/
test_input[24136:24143] = '{32'hc2908cd3, 32'hc1d67087, 32'hc1addf26, 32'hc258897a, 32'h412f285d, 32'h41eadc70, 32'h42c72bb3, 32'hc2abdd10};
test_label[3017] = '{32'hc1addf26};
test_output[3017] = '{32'h42f2a37d};
/*############ DEBUG ############
test_input[24136:24143] = '{-72.2750505385, -26.8049449931, -21.7339594821, -54.1342541329, 10.9473539674, 29.3576355056, 99.5853530627, -85.9317657353};
test_label[3017] = '{-21.7339594821};
test_output[3017] = '{121.319312545};
############ END DEBUG ############*/
test_input[24144:24151] = '{32'hc1c242ac, 32'h42b5eacc, 32'h423a2d75, 32'h4140bd9e, 32'hbff1232e, 32'h42b141f4, 32'h428c43e7, 32'hc2369379};
test_label[3018] = '{32'h42b5eacc};
test_output[3018] = '{32'h3dbe3235};
/*############ DEBUG ############
test_input[24144:24151] = '{-24.2825545343, 90.9585877169, 46.5443900318, 12.0462931725, -1.88388609572, 88.6288184477, 70.1326248561, -45.6440173348};
test_label[3018] = '{90.9585877169};
test_output[3018] = '{0.0928692027706};
############ END DEBUG ############*/
test_input[24152:24159] = '{32'h4247d43f, 32'hc2ad5b8e, 32'hc2bb825a, 32'h428b4b49, 32'hc2895a19, 32'hc118dbcd, 32'hc2ba9c44, 32'h4232aa1d};
test_label[3019] = '{32'hc118dbcd};
test_output[3019] = '{32'h429e66c2};
/*############ DEBUG ############
test_input[24152:24159] = '{49.9572698159, -86.6788165503, -93.7545904002, 69.6470377801, -68.6759719131, -9.55366211054, -93.30520291, 44.6661265863};
test_label[3019] = '{-9.55366211054};
test_output[3019] = '{79.2006998935};
############ END DEBUG ############*/
test_input[24160:24167] = '{32'hc243cc94, 32'hc26da837, 32'hc1a52e5d, 32'hc1c678ed, 32'hc07bd277, 32'hc22023dc, 32'h42a7fa29, 32'hc102d39a};
test_label[3020] = '{32'hc1c678ed};
test_output[3020] = '{32'h42d99864};
/*############ DEBUG ############
test_input[24160:24167] = '{-48.9497848838, -59.4142712183, -20.6476383054, -24.8090449119, -3.93472077414, -40.035019254, 83.9885940667, -8.17666062388};
test_label[3020] = '{-24.8090449119};
test_output[3020] = '{108.797638979};
############ END DEBUG ############*/
test_input[24168:24175] = '{32'h429864e7, 32'hc1f6e9e9, 32'h4290cd35, 32'hc282acf3, 32'hc26f0937, 32'h426e64d4, 32'h428569f9, 32'hc1d92a15};
test_label[3021] = '{32'h4290cd35};
test_output[3021] = '{32'h4074632f};
/*############ DEBUG ############
test_input[24168:24175] = '{76.1970720592, -30.8642135195, 72.4007982712, -65.337793248, -59.7589978469, 59.5984639273, 66.7069813214, -27.1455475963};
test_label[3021] = '{72.4007982712};
test_output[3021] = '{3.81855368223};
############ END DEBUG ############*/
test_input[24176:24183] = '{32'h42c66cdf, 32'h419f9f60, 32'h425a976d, 32'h427f3cb3, 32'h42b52fda, 32'h423c1321, 32'h429ab592, 32'hc1904dbf};
test_label[3022] = '{32'h42b52fda};
test_output[3022] = '{32'h4109e8e9};
/*############ DEBUG ############
test_input[24176:24183] = '{99.2126408369, 19.9528193317, 54.6478775781, 63.8092767148, 90.5934581266, 47.018679166, 77.3546328253, -18.0379627902};
test_label[3022] = '{90.5934581266};
test_output[3022] = '{8.61936330211};
############ END DEBUG ############*/
test_input[24184:24191] = '{32'h4293700b, 32'hc1bd5cc7, 32'hc1a9ab61, 32'hc1225b4a, 32'hc23df502, 32'hc2934204, 32'hc297bd71, 32'hc263297a};
test_label[3023] = '{32'hc1a9ab61};
test_output[3023] = '{32'h42bddae4};
/*############ DEBUG ############
test_input[24184:24191] = '{73.7188372135, -23.6703011768, -21.2086814068, -10.1472872383, -47.4892644939, -73.6289402884, -75.8700036481, -56.790505418};
test_label[3023] = '{-21.2086814068};
test_output[3023] = '{94.9275186203};
############ END DEBUG ############*/
test_input[24192:24199] = '{32'hc23f3645, 32'hc20d5c35, 32'h41e780cc, 32'hc220e039, 32'h42302164, 32'h410c647c, 32'hc1682f4f, 32'h4189df7d};
test_label[3024] = '{32'hc220e039};
test_output[3024] = '{32'h42a880ce};
/*############ DEBUG ############
test_input[24192:24199] = '{-47.8029975846, -35.3400475187, 28.9378889812, -40.2189678262, 44.0326067261, 8.77453198267, -14.5115499779, 17.2341251371};
test_label[3024] = '{-40.2189678262};
test_output[3024] = '{84.2515748305};
############ END DEBUG ############*/
test_input[24200:24207] = '{32'hc28fe417, 32'hc2a4d7ad, 32'hc0b07731, 32'h42c1840c, 32'h4222031b, 32'hc0f4a1d6, 32'hc2193b71, 32'hc1a7ed93};
test_label[3025] = '{32'h4222031b};
test_output[3025] = '{32'h426104fe};
/*############ DEBUG ############
test_input[24200:24207] = '{-71.9454916778, -82.4212427588, -5.51454962891, 96.7579060157, 40.503032624, -7.64475547335, -38.3080481838, -20.9910022395};
test_label[3025] = '{40.503032624};
test_output[3025] = '{56.2548733917};
############ END DEBUG ############*/
test_input[24208:24215] = '{32'hc01480ab, 32'hc0ff0f60, 32'h42c02aa7, 32'hc2aa7d85, 32'hc1de9734, 32'hc2aeeb56, 32'hc0d5f50f, 32'hc1165b7c};
test_label[3026] = '{32'hc2aa7d85};
test_output[3026] = '{32'h43355416};
/*############ DEBUG ############
test_input[24208:24215] = '{-2.32035333141, -7.97062690364, 96.0833052283, -85.2451581683, -27.8238287848, -87.4596368695, -6.68616432218, -9.3973348033};
test_label[3026] = '{-85.2451581683};
test_output[3026] = '{181.328463397};
############ END DEBUG ############*/
test_input[24216:24223] = '{32'hc272a203, 32'h42c6936f, 32'hc2405084, 32'h42a7b4c7, 32'h42a9fe52, 32'h42c14a25, 32'hc1b76722, 32'hc29ab496};
test_label[3027] = '{32'h42a7b4c7};
test_output[3027] = '{32'h41780ebb};
/*############ DEBUG ############
test_input[24216:24223] = '{-60.6582133249, 99.2879541388, -48.0786266793, 83.8530799923, 84.9967226714, 96.6448125101, -22.9253577024, -77.3527045299};
test_label[3027] = '{83.8530799923};
test_output[3027] = '{15.5035960148};
############ END DEBUG ############*/
test_input[24224:24231] = '{32'hc25bc1a5, 32'hc013226d, 32'hc1ba799a, 32'hc21d039f, 32'h3f150626, 32'hbfa2ed73, 32'h418b9742, 32'hc20672b2};
test_label[3028] = '{32'h3f150626};
test_output[3028] = '{32'h4186ef11};
/*############ DEBUG ############
test_input[24224:24231] = '{-54.9391055201, -2.29897619998, -23.3093764971, -39.2535343915, 0.582125096832, -1.27287140233, 17.4488563198, -33.6120083023};
test_label[3028] = '{0.582125096832};
test_output[3028] = '{16.8667312803};
############ END DEBUG ############*/
test_input[24232:24239] = '{32'h411e71a3, 32'h4201d9a0, 32'hc28a8df5, 32'h42157ce8, 32'hc2722982, 32'hc18b2d51, 32'h42b31d7c, 32'hc24641d7};
test_label[3029] = '{32'h42157ce8};
test_output[3029] = '{32'h4250be0f};
/*############ DEBUG ############
test_input[24232:24239] = '{9.90274333017, 32.4625234622, -69.277260949, 37.3719796441, -60.5405352312, -17.397127629, 89.5575836186, -49.5642967451};
test_label[3029] = '{37.3719796441};
test_output[3029] = '{52.1856039744};
############ END DEBUG ############*/
test_input[24240:24247] = '{32'h41764cf6, 32'hc23c149e, 32'h418f2921, 32'hc2a5642e, 32'h42c7005a, 32'h429b9b86, 32'hc29efb09, 32'hc15128f2};
test_label[3030] = '{32'h42c7005a};
test_output[3030] = '{32'h2fcfa3ec};
/*############ DEBUG ############
test_input[24240:24247] = '{15.3937892172, -47.0201339702, 17.8950824381, -82.6956666892, 99.5006886995, 77.8037560987, -79.4902998665, -13.0724965154};
test_label[3030] = '{99.5006886995};
test_output[3030] = '{3.7769554158e-10};
############ END DEBUG ############*/
test_input[24248:24255] = '{32'h4234bdfd, 32'h424e4e1b, 32'hc271935a, 32'hc1d2d65b, 32'hc1332962, 32'hc2b309cf, 32'h4288c977, 32'hc2bcb6fa};
test_label[3031] = '{32'h4288c977};
test_output[3031] = '{32'h3355d40e};
/*############ DEBUG ############
test_input[24248:24255] = '{45.1855369537, 51.5762756496, -60.3938980586, -26.354666404, -11.1976030922, -89.5191560749, 68.393487449, -94.3573735253};
test_label[3031] = '{68.393487449};
test_output[3031] = '{4.97857911744e-08};
############ END DEBUG ############*/
test_input[24256:24263] = '{32'hc211e5d5, 32'hc28ae081, 32'h41e482ba, 32'hc29dfac6, 32'hc1098435, 32'h418d53e3, 32'h4224c8ef, 32'hc2759768};
test_label[3032] = '{32'hc211e5d5};
test_output[3032] = '{32'h429b5762};
/*############ DEBUG ############
test_input[24256:24263] = '{-36.4744435455, -69.438486851, 28.5638306841, -78.9897925813, -8.59477711733, 17.6659609006, 41.1962230603, -61.3978589412};
test_label[3032] = '{-36.4744435455};
test_output[3032] = '{77.6706698703};
############ END DEBUG ############*/
test_input[24264:24271] = '{32'hc29edcb3, 32'hc19b8958, 32'h40ac83b7, 32'h4178fa1c, 32'hc222f349, 32'h424540b1, 32'h4283dde8, 32'h41e6c681};
test_label[3033] = '{32'h4178fa1c};
test_output[3033] = '{32'h42497d48};
/*############ DEBUG ############
test_input[24264:24271] = '{-79.4310515508, -19.4420628424, 5.39107867606, 15.5610618067, -40.7375824048, 49.3131755875, 65.9334070578, 28.8469262815};
test_label[3033] = '{15.5610618067};
test_output[3033] = '{50.3723453117};
############ END DEBUG ############*/
test_input[24272:24279] = '{32'h423709f5, 32'hc2bd51e7, 32'hc2426c0b, 32'hc288d6e6, 32'hbfda5186, 32'h420b1ff9, 32'h4136fdaf, 32'h42823cba};
test_label[3034] = '{32'hc2bd51e7};
test_output[3034] = '{32'h431fc751};
/*############ DEBUG ############
test_input[24272:24279] = '{45.7597250607, -94.6599691736, -48.6055117813, -68.4197198163, -1.70561292009, 34.7812245886, 11.4369348312, 65.118607783};
test_label[3034] = '{-94.6599691736};
test_output[3034] = '{159.778576961};
############ END DEBUG ############*/
test_input[24280:24287] = '{32'h42a33dd8, 32'h4233d382, 32'hc226506a, 32'h4284c7fc, 32'h4221d115, 32'h40bd1d64, 32'hc22c86b5, 32'hc25e940d};
test_label[3035] = '{32'hc22c86b5};
test_output[3035] = '{32'h42f98133};
/*############ DEBUG ############
test_input[24280:24287] = '{81.6207899573, 44.9565496358, -41.5785295972, 66.390593265, 40.4541803892, 5.9098378232, -43.1315515348, -55.6445796492};
test_label[3035] = '{-43.1315515348};
test_output[3035] = '{124.752341735};
############ END DEBUG ############*/
test_input[24288:24295] = '{32'h4205cb2f, 32'hc260ac07, 32'h40b5ccc9, 32'h42b542a3, 32'h4137718c, 32'h42a15b28, 32'hc2baf16c, 32'hc2aeb7b8};
test_label[3036] = '{32'h4205cb2f};
test_output[3036] = '{32'h4264ba24};
/*############ DEBUG ############
test_input[24288:24295] = '{33.4484230084, -56.1679954657, 5.6812480258, 90.6301532882, 11.4652209347, 80.6780422914, -93.4715244267, -87.3588220257};
test_label[3036] = '{33.4484230084};
test_output[3036] = '{57.1817779057};
############ END DEBUG ############*/
test_input[24296:24303] = '{32'h41782a10, 32'h421dacd2, 32'hc208225c, 32'h42bcbe7d, 32'h42639109, 32'h4215d6fb, 32'hc09b25e3, 32'h42bfe068};
test_label[3037] = '{32'h4215d6fb};
test_output[3037] = '{32'h426aac08};
/*############ DEBUG ############
test_input[24296:24303] = '{15.5102693005, 39.418770986, -34.0335533864, 94.3720474627, 56.8916364053, 37.45994326, -4.84837495947, 95.938292671};
test_label[3037] = '{37.45994326};
test_output[3037] = '{58.6680005548};
############ END DEBUG ############*/
test_input[24304:24311] = '{32'hc2aeb116, 32'hc00cb02b, 32'h41877821, 32'hc2c72a23, 32'h427a8fd6, 32'hc1aac4a6, 32'h4000acd2, 32'hc268021b};
test_label[3038] = '{32'hc00cb02b};
test_output[3038] = '{32'h4281ad6c};
/*############ DEBUG ############
test_input[24304:24311] = '{-87.3458746969, -2.19825245789, 16.9336565848, -99.5822955846, 62.6404645206, -21.3460205539, 2.01054804934, -58.0020544455};
test_label[3038] = '{-2.19825245789};
test_output[3038] = '{64.8387169785};
############ END DEBUG ############*/
test_input[24312:24319] = '{32'h40544a08, 32'h421a8c32, 32'h41c9de54, 32'h4297c0f0, 32'hc166644b, 32'h40c05825, 32'h42c49bb2, 32'h428bd7d7};
test_label[3039] = '{32'h428bd7d7};
test_output[3039] = '{32'h41e30f6b};
/*############ DEBUG ############
test_input[24312:24319] = '{3.31701849498, 38.6369087858, 25.2335587512, 75.8768296586, -14.3994851345, 6.01076001427, 98.3040940359, 69.9215659711};
test_label[3039] = '{69.9215659711};
test_output[3039] = '{28.3825280649};
############ END DEBUG ############*/
test_input[24320:24327] = '{32'hc1071d03, 32'hc2a80017, 32'h421e5c4c, 32'h4290215f, 32'h41672ff3, 32'hbe393d38, 32'hc29e1f5e, 32'hc28fb11f};
test_label[3040] = '{32'hbe393d38};
test_output[3040] = '{32'h42907dfe};
/*############ DEBUG ############
test_input[24320:24327] = '{-8.44458295097, -84.0001792113, 39.5901320758, 72.0651797239, 14.4492062545, -0.180897589123, -79.0612671405, -71.845939404};
test_label[3040] = '{-0.180897589123};
test_output[3040] = '{72.246077313};
############ END DEBUG ############*/
test_input[24328:24335] = '{32'h42509c92, 32'h412359c8, 32'hc2284346, 32'h41e1af66, 32'h4255dfd8, 32'hc2782a03, 32'hc1c887f3, 32'hc14c7350};
test_label[3041] = '{32'h41e1af66};
test_output[3041] = '{32'h41cbf708};
/*############ DEBUG ############
test_input[24328:24335] = '{52.1528990778, 10.2094192397, -42.0656967373, 28.2106428659, 53.4685955854, -62.0410264256, -25.0663823531, -12.7781526447};
test_label[3041] = '{28.2106428659};
test_output[3041] = '{25.4956202012};
############ END DEBUG ############*/
test_input[24336:24343] = '{32'h4286e95b, 32'h4293b2af, 32'h426a8348, 32'hc2b7c385, 32'h42b6a1cc, 32'hc186cef7, 32'h423d6a42, 32'h41db7a82};
test_label[3042] = '{32'h426a8348};
test_output[3042] = '{32'h4202c051};
/*############ DEBUG ############
test_input[24336:24343] = '{67.4557758338, 73.8489946116, 58.6282034896, -91.8818709786, 91.3160105503, -16.8510567688, 47.3537666459, 27.4348187103};
test_label[3042] = '{58.6282034896};
test_output[3042] = '{32.6878070868};
############ END DEBUG ############*/
test_input[24344:24351] = '{32'hc28a9c38, 32'hc28fecd0, 32'hc291a917, 32'hc1ab6e8a, 32'h426d18e5, 32'h4262d4c3, 32'hc0dec0f1, 32'hc26fcbbf};
test_label[3043] = '{32'h4262d4c3};
test_output[3043] = '{32'h4028fe81};
/*############ DEBUG ############
test_input[24344:24351] = '{-69.3051171713, -71.9625235772, -72.8302516144, -21.4289735099, 59.2743128244, 56.7077735381, -6.96105245805, -59.9489709317};
test_label[3043] = '{56.7077735381};
test_output[3043] = '{2.64053377586};
############ END DEBUG ############*/
test_input[24352:24359] = '{32'hc226b848, 32'hc25e7dbd, 32'h4156cef9, 32'h4222097a, 32'h42915d9f, 32'h42446fe1, 32'hc2b4c119, 32'h4212a1c1};
test_label[3044] = '{32'h42915d9f};
test_output[3044] = '{32'h2e7e5d60};
/*############ DEBUG ############
test_input[24352:24359] = '{-41.6799631266, -55.6227907068, 13.4255308349, 40.5092546729, 72.682857357, 49.1092560953, -90.3771431878, 36.6579615758};
test_label[3044] = '{72.682857357};
test_output[3044] = '{5.78358472242e-11};
############ END DEBUG ############*/
test_input[24360:24367] = '{32'h414417c7, 32'hc1fede1d, 32'h426dffd3, 32'h419c3921, 32'hc2c6c996, 32'h42c65280, 32'hc2c597bd, 32'h428b5993};
test_label[3045] = '{32'hc1fede1d};
test_output[3045] = '{32'h43030504};
/*############ DEBUG ############
test_input[24360:24367] = '{12.2558047516, -31.8584530578, 59.4998273796, 19.5278946109, -99.3937192289, 99.1611324068, -98.7963623735, 69.6749487754};
test_label[3045] = '{-31.8584530578};
test_output[3045] = '{131.019585465};
############ END DEBUG ############*/
test_input[24368:24375] = '{32'hc276554e, 32'hc28348f7, 32'hc07f8678, 32'hc2bbf6cd, 32'hc0c951de, 32'h42bbafce, 32'hc264db2d, 32'h425c6761};
test_label[3046] = '{32'hc2bbf6cd};
test_output[3046] = '{32'h433bd34e};
/*############ DEBUG ############
test_input[24368:24375] = '{-61.5833036363, -65.6425098488, -3.99258233512, -93.9820355463, -6.29124348233, 93.8433664185, -57.2140370532, 55.1009549256};
test_label[3046] = '{-93.9820355463};
test_output[3046] = '{187.825401965};
############ END DEBUG ############*/
test_input[24376:24383] = '{32'hc1f702ea, 32'h41c74b7f, 32'h421bcdd6, 32'hc2207432, 32'h40a1e1fa, 32'hc2c06600, 32'hc2b20fe7, 32'hc21e3b43};
test_label[3047] = '{32'h40a1e1fa};
test_output[3047] = '{32'h42079197};
/*############ DEBUG ############
test_input[24376:24383] = '{-30.8764220005, 24.9118624422, 38.9510117956, -40.1134718156, 5.05883493809, -96.1992180973, -89.031057369, -39.5578740291};
test_label[3047] = '{5.05883493809};
test_output[3047] = '{33.8921776571};
############ END DEBUG ############*/
test_input[24384:24391] = '{32'hc1b01a16, 32'hc12bf33a, 32'hc2567660, 32'h4151093c, 32'hc210ee06, 32'hc1b16810, 32'hc1b85935, 32'hc2212ee8};
test_label[3048] = '{32'h4151093c};
test_output[3048] = '{32'h2e4873c0};
/*############ DEBUG ############
test_input[24384:24391] = '{-22.0127370073, -10.7468819452, -53.6156001934, 13.0647543526, -36.232443037, -22.1758116991, -23.0435578542, -40.2958070057};
test_label[3048] = '{13.0647543526};
test_output[3048] = '{4.55775417418e-11};
############ END DEBUG ############*/
test_input[24392:24399] = '{32'hc10fd45d, 32'hc21cef81, 32'hc16ac1ce, 32'h42947b4d, 32'h42bf1902, 32'hc2201879, 32'h4219d6c0, 32'h4274ef76};
test_label[3049] = '{32'h4219d6c0};
test_output[3049] = '{32'h42645b44};
/*############ DEBUG ############
test_input[24392:24399] = '{-8.98934691842, -39.2338914926, -14.6723156279, 74.2408221493, 95.5488469934, -40.0238986073, 38.4597185271, 61.2338500542};
test_label[3049] = '{38.4597185271};
test_output[3049] = '{57.0891284668};
############ END DEBUG ############*/
test_input[24400:24407] = '{32'hc2604d55, 32'h429e8aae, 32'h418177fa, 32'hc2b74a38, 32'h41aacd07, 32'hc2c79943, 32'h415ad480, 32'h4209a56e};
test_label[3050] = '{32'h415ad480};
test_output[3050] = '{32'h4283301e};
/*############ DEBUG ############
test_input[24400:24407] = '{-56.0755195271, 79.2708564982, 16.183583256, -91.6449607023, 21.3501106494, -99.7993370083, 13.6768797699, 34.4115515624};
test_label[3050] = '{13.6768797699};
test_output[3050] = '{65.5939767282};
############ END DEBUG ############*/
test_input[24408:24415] = '{32'h42b44026, 32'h41220540, 32'h428c97db, 32'hc1fde198, 32'hc022b153, 32'h4103fe90, 32'h42bd52ee, 32'hc22bf05c};
test_label[3051] = '{32'hc22bf05c};
test_output[3051] = '{32'h4309a848};
/*############ DEBUG ############
test_input[24408:24415] = '{90.1252881872, 10.1262814552, 70.2965914053, -31.7351524296, -2.54207310959, 8.24964903166, 94.6619686589, -42.9847249825};
test_label[3051] = '{-42.9847249825};
test_output[3051] = '{137.657345603};
############ END DEBUG ############*/
test_input[24416:24423] = '{32'h42299265, 32'h4220974b, 32'h420e7868, 32'hc297d33b, 32'h427f7dc7, 32'hc126224d, 32'hc2a35149, 32'h4281b45d};
test_label[3052] = '{32'h4220974b};
test_output[3052] = '{32'h41c82fd5};
/*############ DEBUG ############
test_input[24416:24423] = '{42.3929628141, 40.1477489352, 35.6175853322, -75.9125570771, 63.872830969, -10.3833737604, -81.6587581055, 64.8522706897};
test_label[3052] = '{40.1477489352};
test_output[3052] = '{25.0233546406};
############ END DEBUG ############*/
test_input[24424:24431] = '{32'hc212dae6, 32'h4213f64b, 32'hc283fc66, 32'h422c7c0d, 32'hc285ca09, 32'hc22f39ad, 32'hc298a03e, 32'hc0a91582};
test_label[3053] = '{32'hc285ca09};
test_output[3053] = '{32'h42dc092c};
/*############ DEBUG ############
test_input[24424:24431] = '{-36.7137675326, 36.9905190211, -65.9929647958, 43.1211437226, -66.894596812, -43.8063251927, -76.3129704548, -5.28387558047};
test_label[3053] = '{-66.894596812};
test_output[3053] = '{110.017913394};
############ END DEBUG ############*/
test_input[24432:24439] = '{32'hc2c38359, 32'h429d34e9, 32'hc2b3516e, 32'hc22e4a78, 32'h42859d08, 32'hc163032f, 32'h42ba0c8c, 32'h42c5d27b};
test_label[3054] = '{32'hc2b3516e};
test_output[3054] = '{32'h433c92aa};
/*############ DEBUG ############
test_input[24432:24439] = '{-97.7565349328, 78.6033421587, -89.6590457441, -43.5727250832, 66.8067040583, -14.188276808, 93.0245074614, 98.9110936489};
test_label[3054] = '{-89.6590457441};
test_output[3054] = '{188.572911986};
############ END DEBUG ############*/
test_input[24440:24447] = '{32'h42bab193, 32'hc2aad9b4, 32'hc2971b36, 32'hc2b38328, 32'h42b42051, 32'hc293bf3b, 32'h411a6ba1, 32'hc2a515c1};
test_label[3055] = '{32'hc2aad9b4};
test_output[3055] = '{32'h4332cf10};
/*############ DEBUG ############
test_input[24440:24447] = '{93.3468275558, -85.425201235, -75.5531440945, -89.7561627228, 90.0631198496, -73.8734942617, 9.65127622466, -82.5424875861};
test_label[3055] = '{-85.425201235};
test_output[3055] = '{178.808832162};
############ END DEBUG ############*/
test_input[24448:24455] = '{32'h417fd436, 32'hc1b4a35c, 32'hc2a6112b, 32'h42426e41, 32'h40365aa5, 32'hc28e983c, 32'hc1a9ccaf, 32'h419f5762};
test_label[3056] = '{32'h417fd436};
test_output[3056] = '{32'h42027934};
/*############ DEBUG ############
test_input[24448:24455] = '{15.9893097591, -22.579765624, -83.0335342498, 48.6076713003, 2.84928245227, -71.2973315475, -21.2249440624, 19.9176672909};
test_label[3056] = '{15.9893097591};
test_output[3056] = '{32.6183615411};
############ END DEBUG ############*/
test_input[24456:24463] = '{32'hc29873b8, 32'h40818620, 32'h40c55e84, 32'hc2bb38c9, 32'hc2978232, 32'h41a41fb9, 32'h42c4164c, 32'hc22d2dc3};
test_label[3057] = '{32'hc22d2dc3};
test_output[3057] = '{32'h430d5697};
/*############ DEBUG ############
test_input[24456:24463] = '{-76.2260114287, 4.04762285441, 6.16778778551, -93.6109103473, -75.7542876999, 20.5154887301, 98.0435468029, -43.2946902817};
test_label[3057] = '{-43.2946902817};
test_output[3057] = '{141.338237085};
############ END DEBUG ############*/
test_input[24464:24471] = '{32'h42aab322, 32'h42a87fd5, 32'h42b58c71, 32'hc21eb296, 32'h427f6d75, 32'hc2c5ee2b, 32'hc2899513, 32'h428684d2};
test_label[3058] = '{32'hc21eb296};
test_output[3058] = '{32'h4302745e};
/*############ DEBUG ############
test_input[24464:24471] = '{85.3498692008, 84.2496693562, 90.7743030637, -39.6744015658, 63.85689066, -98.9651747217, -68.7911570224, 67.2594181392};
test_label[3058] = '{-39.6744015658};
test_output[3058] = '{130.45456186};
############ END DEBUG ############*/
test_input[24472:24479] = '{32'hc1fe5d76, 32'h4232592a, 32'h42bd1983, 32'h411a09d1, 32'h41ceb822, 32'hc28e9b31, 32'h42ba80b8, 32'h42bc170b};
test_label[3059] = '{32'hc28e9b31};
test_output[3059] = '{32'h43267b7e};
/*############ DEBUG ############
test_input[24472:24479] = '{-31.795634815, 44.5870755656, 94.5498287129, 9.62739667204, 25.8399077549, -71.3031100411, 93.2514012299, 94.0450075617};
test_label[3059] = '{-71.3031100411};
test_output[3059] = '{166.482386641};
############ END DEBUG ############*/
test_input[24480:24487] = '{32'h41aa1862, 32'h42963063, 32'hc29391f4, 32'hc1263270, 32'h418ef4bb, 32'h41cbc72e, 32'hc2aea548, 32'hc17b356a};
test_label[3060] = '{32'h418ef4bb};
test_output[3060] = '{32'h4264e669};
/*############ DEBUG ############
test_input[24480:24487] = '{21.261905555, 75.094507529, -73.7850665321, -10.3873134519, 17.8694967292, 25.4722553555, -87.3228184752, -15.7005410132};
test_label[3060] = '{17.8694967292};
test_output[3060] = '{57.2250107999};
############ END DEBUG ############*/
test_input[24488:24495] = '{32'hc2400e2f, 32'hc2141a30, 32'h41ce1e27, 32'hc29ad844, 32'hc118738c, 32'h4264c399, 32'h42bfd6ef, 32'hc191330f};
test_label[3061] = '{32'hc29ad844};
test_output[3061] = '{32'h432d579a};
/*############ DEBUG ############
test_input[24488:24495] = '{-48.0138502324, -37.0255748191, 25.764723265, -77.4223949769, -9.52820972748, 57.1910140586, 95.9197917084, -18.1499304001};
test_label[3061] = '{-77.4223949769};
test_output[3061] = '{173.342186685};
############ END DEBUG ############*/
test_input[24496:24503] = '{32'hc2756bc4, 32'h42ab166e, 32'h42a3c86d, 32'hc2bc77c9, 32'hc241c67d, 32'h403cd247, 32'h41e4ba28, 32'hc2aab74d};
test_label[3062] = '{32'h42ab166e};
test_output[3062] = '{32'h3cd1b623};
/*############ DEBUG ############
test_input[24496:24503] = '{-61.3552416025, 85.543806475, 81.8914528101, -94.2339520354, -48.4438353279, 2.95033432841, 28.5908959507, -85.3580106235};
test_label[3062] = '{85.543806475};
test_output[3062] = '{0.0255995439404};
############ END DEBUG ############*/
test_input[24504:24511] = '{32'hc1369a38, 32'h428ee217, 32'hc299c2b9, 32'hc28789e7, 32'hc2ac7d71, 32'hc1b427f2, 32'h40fe4b42, 32'h42bd41ad};
test_label[3063] = '{32'hc2ac7d71};
test_output[3063] = '{32'h4334df8f};
/*############ DEBUG ############
test_input[24504:24511] = '{-11.412650858, 71.4415790067, -76.8803172699, -67.7693408241, -86.2449997057, -22.5195035976, 7.94668666255, 94.6282767823};
test_label[3063] = '{-86.2449997057};
test_output[3063] = '{180.873276488};
############ END DEBUG ############*/
test_input[24512:24519] = '{32'hc2b3e68c, 32'hc1a4fa58, 32'hc14379b3, 32'hc10a6e67, 32'h42a71fff, 32'hc2b925c0, 32'hc1f6c642, 32'hc2c15594};
test_label[3064] = '{32'hc2c15594};
test_output[3064] = '{32'h43343aca};
/*############ DEBUG ############
test_input[24512:24519] = '{-89.950284236, -20.6222384523, -12.217211683, -8.65195351942, 83.5624927819, -92.5737280622, -30.846805763, -96.6671479599};
test_label[3064] = '{-96.6671479599};
test_output[3064] = '{180.229640742};
############ END DEBUG ############*/
test_input[24520:24527] = '{32'hc290e64e, 32'hc18fd18a, 32'h41e88da1, 32'h429206a5, 32'h42a2222f, 32'h420822ae, 32'hc238b3a3, 32'hc2c62e67};
test_label[3065] = '{32'h420822ae};
test_output[3065] = '{32'h423c2203};
/*############ DEBUG ############
test_input[24520:24527] = '{-72.4498168127, -17.977313361, 29.0691541062, 73.012976926, 81.0667634552, 34.0338668228, -46.1754277856, -99.0906269128};
test_label[3065] = '{34.0338668228};
test_output[3065] = '{47.0332144778};
############ END DEBUG ############*/
test_input[24528:24535] = '{32'h42c6b155, 32'hc1dea530, 32'hc1fc628c, 32'hc20c6381, 32'hc1400a36, 32'h4275ac72, 32'h42076cd5, 32'hc2a29687};
test_label[3066] = '{32'h42c6b155};
test_output[3066] = '{32'h80000000};
/*############ DEBUG ############
test_input[24528:24535] = '{99.3463533184, -27.830658786, -31.5481187319, -35.0971699196, -12.0024930295, 61.4184040789, 33.8562800183, -81.29399496};
test_label[3066] = '{99.3463533184};
test_output[3066] = '{-0.0};
############ END DEBUG ############*/
test_input[24536:24543] = '{32'hc0d9e1ae, 32'h41b0faaf, 32'hc2798f4c, 32'hc250b5ac, 32'hc2886e10, 32'h428df794, 32'h42972255, 32'h41560431};
test_label[3067] = '{32'h428df794};
test_output[3067] = '{32'h4092ff54};
/*############ DEBUG ############
test_input[24536:24543] = '{-6.8087986016, 22.1224044593, -62.3899390506, -52.1774146954, -68.2149645476, 70.9835507896, 75.5670515713, 13.3760236397};
test_label[3067] = '{70.9835507896};
test_output[3067] = '{4.59366797902};
############ END DEBUG ############*/
test_input[24544:24551] = '{32'h41e3a418, 32'h41060b69, 32'h4291091b, 32'h420b9579, 32'h411a6099, 32'h42a420bb, 32'h41777195, 32'h41427c0f};
test_label[3068] = '{32'h41777195};
test_output[3068] = '{32'h42853292};
/*############ DEBUG ############
test_input[24544:24551] = '{28.4551245237, 8.37778542206, 72.5177821349, 34.8959682251, 9.64858304406, 82.0639304856, 15.4652302307, 12.1552880282};
test_label[3068] = '{15.4652302307};
test_output[3068] = '{66.5987717284};
############ END DEBUG ############*/
test_input[24552:24559] = '{32'h42be895d, 32'h4187206b, 32'hc1a5d867, 32'h41ed9fdd, 32'hc1d21f61, 32'h41eefed0, 32'h3f862c7f, 32'h41649ddc};
test_label[3069] = '{32'h41eefed0};
test_output[3069] = '{32'h4282c9a9};
/*############ DEBUG ############
test_input[24552:24559] = '{95.2682893091, 16.8908297176, -20.7306659567, 29.7030578175, -26.2653210069, 29.8744192874, 1.04823293081, 14.2885397553};
test_label[3069] = '{29.8744192874};
test_output[3069] = '{65.3938700217};
############ END DEBUG ############*/
test_input[24560:24567] = '{32'hc2398242, 32'hc27818db, 32'h42a471ac, 32'h41888c74, 32'hc28a4368, 32'h42ab81c5, 32'hc111aca6, 32'h4195d310};
test_label[3070] = '{32'hc28a4368};
test_output[3070] = '{32'h431ae9f9};
/*############ DEBUG ############
test_input[24560:24567] = '{-46.3772048791, -62.0242711761, 82.222017663, 17.0685801387, -69.1316563948, 85.7534593609, -9.10465006584, 18.7280572216};
test_label[3070] = '{-69.1316563948};
test_output[3070] = '{154.913958474};
############ END DEBUG ############*/
test_input[24568:24575] = '{32'h41f8a4ff, 32'h4291baac, 32'hc2535910, 32'h42aea807, 32'hc2a5c581, 32'h41f61755, 32'h41c48654, 32'h417f283c};
test_label[3071] = '{32'h41f8a4ff};
test_output[3071] = '{32'h4260fd8e};
/*############ DEBUG ############
test_input[24568:24575] = '{31.0805636237, 72.8645966605, -52.8369737728, 87.3281753618, -82.8857494304, 30.7613920644, 24.5655899012, 15.9473230116};
test_label[3071] = '{31.0805636237};
test_output[3071] = '{56.2476122611};
############ END DEBUG ############*/
test_input[24576:24583] = '{32'h42088b28, 32'h426daf0f, 32'h429a8ed3, 32'h42b5653b, 32'hc1a32061, 32'hc1d9eb70, 32'hc178cfc1, 32'h420442c9};
test_label[3072] = '{32'hc1d9eb70};
test_output[3072] = '{32'h42ebe017};
/*############ DEBUG ############
test_input[24576:24583] = '{34.1358943187, 59.420956057, 77.2789562947, 90.6977156025, -20.3908091678, -27.2399590394, -15.5507212887, 33.0652202178};
test_label[3072] = '{-27.2399590394};
test_output[3072] = '{117.937676129};
############ END DEBUG ############*/
test_input[24584:24591] = '{32'hc269fbe4, 32'hc285059f, 32'hc2c6366d, 32'hc28f2fc9, 32'h41e5705f, 32'h42c38556, 32'h40a43a87, 32'h4245e7b5};
test_label[3073] = '{32'h42c38556};
test_output[3073] = '{32'h80000000};
/*############ DEBUG ############
test_input[24584:24591] = '{-58.4959885099, -66.5109814656, -99.1063007716, -71.5933332676, 28.6798691559, 97.7604231525, 5.13214444425, 49.4762779452};
test_label[3073] = '{97.7604231525};
test_output[3073] = '{-0.0};
############ END DEBUG ############*/
test_input[24592:24599] = '{32'h41e00c19, 32'hc1d291dc, 32'hc15389b7, 32'hc2852254, 32'hc22ca62a, 32'h4060d5a0, 32'h41caccfd, 32'hc1b71bf1};
test_label[3074] = '{32'hc1b71bf1};
test_output[3074] = '{32'h424bd988};
/*############ DEBUG ############
test_input[24592:24599] = '{28.0059061118, -26.3212201551, -13.2211221335, -66.5670507648, -43.1622712927, 3.51303860699, 25.3500920249, -22.8886428602};
test_label[3074] = '{-22.8886428602};
test_output[3074] = '{50.9624334199};
############ END DEBUG ############*/
test_input[24600:24607] = '{32'hc253a430, 32'h4285a3ae, 32'h41ee29be, 32'hc1973626, 32'hc21b0b3d, 32'hbf88cb33, 32'hc23771df, 32'h426b5750};
test_label[3075] = '{32'h426b5750};
test_output[3075] = '{32'h40ff832d};
/*############ DEBUG ############
test_input[24600:24607] = '{-52.9103390557, 66.8196882119, 29.770382723, -18.9014396494, -38.7609730763, -1.06870113121, -45.8612018947, 58.835266041};
test_label[3075] = '{58.835266041};
test_output[3075] = '{7.98476284218};
############ END DEBUG ############*/
test_input[24608:24615] = '{32'hc23a1ce7, 32'hc286bd22, 32'h420442d6, 32'h40edbd59, 32'hc2c1dddb, 32'h42842beb, 32'h421fa7a0, 32'hc25af094};
test_label[3076] = '{32'h421fa7a0};
test_output[3076] = '{32'h41d1606b};
/*############ DEBUG ############
test_input[24608:24615] = '{-46.5282268131, -67.3693998169, 33.065271188, 7.4293638038, -96.9333138486, 66.0857760885, 39.9136965184, -54.7349403647};
test_label[3076] = '{39.9136965184};
test_output[3076] = '{26.17207957};
############ END DEBUG ############*/
test_input[24616:24623] = '{32'h421d33ee, 32'h424a2823, 32'hc28546e9, 32'h42b6d227, 32'h4189912f, 32'h41f625f9, 32'h42c631b3, 32'h417f7b27};
test_label[3077] = '{32'h42b6d227};
test_output[3077] = '{32'h40f5fc8e};
/*############ DEBUG ############
test_input[24616:24623] = '{39.3007114916, 50.5391974065, -66.638495669, 91.4104507549, 17.1958907093, 30.7685412533, 99.0970715416, 15.9675664976};
test_label[3077] = '{91.4104507549};
test_output[3077] = '{7.68707960776};
############ END DEBUG ############*/
test_input[24624:24631] = '{32'h424eee0f, 32'hc18be1b9, 32'h426dc205, 32'hbfd9d73b, 32'h427fbc11, 32'hc1ddc597, 32'hc26cc87d, 32'h42c0d818};
test_label[3078] = '{32'hc1ddc597};
test_output[3078] = '{32'h42f8497e};
/*############ DEBUG ############
test_input[24624:24631] = '{51.7324777417, -17.4852162274, 59.4394705247, -1.70188084652, 63.9336575428, -27.7214801823, -59.1957899972, 96.422056354};
test_label[3078] = '{-27.7214801823};
test_output[3078] = '{124.143536536};
############ END DEBUG ############*/
test_input[24632:24639] = '{32'hc188b4c1, 32'h427b61db, 32'hc2805002, 32'hc2a30469, 32'h429186fd, 32'h42c35669, 32'hc28d119a, 32'h41871817};
test_label[3079] = '{32'h42c35669};
test_output[3079] = '{32'h2d865300};
/*############ DEBUG ############
test_input[24632:24639] = '{-17.0882596842, 62.8455608335, -64.1562682352, -81.5086135449, 72.7636485956, 97.6687707473, -70.5343794578, 16.8867621686};
test_label[3079] = '{97.6687707473};
test_output[3079] = '{1.52708956592e-11};
############ END DEBUG ############*/
test_input[24640:24647] = '{32'h426a5d09, 32'hc23aaa40, 32'hc2264b1e, 32'hc2a13022, 32'hc21035f4, 32'h3fa28f78, 32'hc2269ea8, 32'h415db358};
test_label[3080] = '{32'hc2a13022};
test_output[3080] = '{32'h430b2f53};
/*############ DEBUG ############
test_input[24640:24647] = '{58.5908533509, -46.6662615588, -41.5733574258, -80.5940088803, -36.0526870393, 1.27000336283, -41.6549372518, 13.8562855287};
test_label[3080] = '{-80.5940088803};
test_output[3080] = '{139.184862231};
############ END DEBUG ############*/
test_input[24648:24655] = '{32'hc06eed23, 32'h41c42a10, 32'h42a2c9fc, 32'hc2aab6b6, 32'hc1e72f73, 32'hc20f0c45, 32'hc200bfb8, 32'h42c0ec4b};
test_label[3081] = '{32'h41c42a10};
test_output[3081] = '{32'h428fe1c7};
/*############ DEBUG ############
test_input[24648:24655] = '{-3.73322368172, 24.5205375244, 81.3944991769, -85.3568597078, -28.8981686737, -35.7619822537, -32.1872254774, 96.4615110249};
test_label[3081] = '{24.5205375244};
test_output[3081] = '{71.9409737866};
############ END DEBUG ############*/
test_input[24656:24663] = '{32'hc1debad2, 32'h4291c405, 32'hc217888c, 32'h41b83745, 32'hc2b7e9f2, 32'hc29c047c, 32'h42043248, 32'hc2584a47};
test_label[3082] = '{32'hc1debad2};
test_output[3082] = '{32'h42c972b9};
/*############ DEBUG ############
test_input[24656:24663] = '{-27.8412205989, 72.8828493376, -37.8833459669, 23.0269870087, -91.9569250673, -78.00875477, 33.0491032856, -54.0725376378};
test_label[3082] = '{-27.8412205989};
test_output[3082] = '{100.724069936};
############ END DEBUG ############*/
test_input[24664:24671] = '{32'hc1d12cf9, 32'hc24dfedd, 32'hc03fc026, 32'hc27a8512, 32'hc18b3eab, 32'h404fc617, 32'h42b86140, 32'h40862478};
test_label[3083] = '{32'hc1d12cf9};
test_output[3083] = '{32'h42ecac7f};
/*############ DEBUG ############
test_input[24664:24671] = '{-26.1469589386, -51.4988895706, -2.99610278395, -62.6299497282, -17.4055990961, 3.24646546774, 92.1899439328, 4.19195159772};
test_label[3083] = '{-26.1469589386};
test_output[3083] = '{118.336902871};
############ END DEBUG ############*/
test_input[24672:24679] = '{32'hc28770c2, 32'hc1bc6c81, 32'hc26dc442, 32'hc276bc7e, 32'hc2aa3fed, 32'h4213fe47, 32'h42a1200e, 32'h42863183};
test_label[3084] = '{32'hc276bc7e};
test_output[3084] = '{32'h430e3f26};
/*############ DEBUG ############
test_input[24672:24679] = '{-67.7202312322, -23.5529809643, -59.4416579663, -61.6840743399, -85.1248587113, 36.9983185636, 80.5626044319, 67.0967037628};
test_label[3084] = '{-61.6840743399};
test_output[3084] = '{142.24668019};
############ END DEBUG ############*/
test_input[24680:24687] = '{32'h41d84b2f, 32'hc20aefcf, 32'hc0c09ded, 32'h42593967, 32'hc29c6f86, 32'h40b66a08, 32'h40da1d0c, 32'hc2203a73};
test_label[3085] = '{32'hc20aefcf};
test_output[3085] = '{32'h42b2149b};
/*############ DEBUG ############
test_input[24680:24687] = '{27.0367116197, -34.7341879584, -6.01927794015, 54.3060559739, -78.2178168388, 5.70044343011, 6.81604590388, -40.0570797685};
test_label[3085] = '{-34.7341879584};
test_output[3085] = '{89.0402439322};
############ END DEBUG ############*/
test_input[24688:24695] = '{32'h421e33aa, 32'h42b281db, 32'h419c65cb, 32'hc2a684ee, 32'h4188fd60, 32'hc2118875, 32'hc2b4c516, 32'h425161a0};
test_label[3086] = '{32'h419c65cb};
test_output[3086] = '{32'h428b6868};
/*############ DEBUG ############
test_input[24688:24695] = '{39.5504529616, 89.2536252079, 19.5497031438, -83.2596308454, 17.1237187851, -36.3832596964, -90.3849369696, 52.3453357262};
test_label[3086] = '{19.5497031438};
test_output[3086] = '{69.703922064};
############ END DEBUG ############*/
test_input[24696:24703] = '{32'hc24bb5f0, 32'hc0c7301a, 32'h42b3476c, 32'hc1d8981f, 32'hc24b2d8e, 32'hc2bd0769, 32'h42847f51, 32'h425b5982};
test_label[3087] = '{32'h42b3476c};
test_output[3087] = '{32'h2e98a910};
/*############ DEBUG ############
test_input[24696:24703] = '{-50.9276725517, -6.22462199845, 89.639496857, -27.0742772461, -50.7944853612, -94.5144732755, 66.2486666715, 54.8374106081};
test_label[3087] = '{89.639496857};
test_output[3087] = '{6.94219126653e-11};
############ END DEBUG ############*/
test_input[24704:24711] = '{32'h42532455, 32'hc2ba1d21, 32'h42b6739d, 32'hc245b8be, 32'h426b2617, 32'hc273f3c5, 32'h41be922c, 32'hc223ae19};
test_label[3088] = '{32'h42b6739d};
test_output[3088] = '{32'h28120000};
/*############ DEBUG ############
test_input[24704:24711] = '{52.7854787729, -93.056890291, 91.2258046273, -49.4304121939, 58.7871960057, -60.9880569365, 23.8213723903, -40.9200169006};
test_label[3088] = '{91.2258046273};
test_output[3088] = '{8.10462807976e-15};
############ END DEBUG ############*/
test_input[24712:24719] = '{32'hc293f48e, 32'h41d80b24, 32'h42837fa2, 32'h4245c074, 32'h41ee9ef1, 32'hc1f525b2, 32'hc2932e9e, 32'hc26e2fd2};
test_label[3089] = '{32'h4245c074};
test_output[3089] = '{32'h41827da2};
/*############ DEBUG ############
test_input[24712:24719] = '{-73.9776486262, 27.005439411, 65.749285566, 49.4379423884, 29.8276079884, -30.643405674, -73.5910510453, -59.5466978279};
test_label[3089] = '{49.4379423884};
test_output[3089] = '{16.31134326};
############ END DEBUG ############*/
test_input[24720:24727] = '{32'hc1cf3d91, 32'hc2b0c55f, 32'h41f91652, 32'h42625ca5, 32'h423fa934, 32'hc2570d5a, 32'hc26b8846, 32'h41e761ec};
test_label[3090] = '{32'h41e761ec};
test_output[3090] = '{32'h41dd57b7};
/*############ DEBUG ############
test_input[24720:24727] = '{-25.9050614396, -88.3854878244, 31.1358981534, 56.5904725979, 47.9152388596, -53.7630393521, -58.8830779809, 28.9228129776};
test_label[3090] = '{28.9228129776};
test_output[3090] = '{27.6678303687};
############ END DEBUG ############*/
test_input[24728:24735] = '{32'hc2be0eea, 32'hc1521e6d, 32'h423800ec, 32'hc263c395, 32'h428ebdd3, 32'hc25eb0a5, 32'hc257542e, 32'h42b91706};
test_label[3091] = '{32'hc257542e};
test_output[3091] = '{32'h4312608e};
/*############ DEBUG ############
test_input[24728:24735] = '{-95.0291260499, -13.1324282868, 46.0009005906, -56.9409989879, 71.370749164, -55.672505142, -53.8322057263, 92.5449673429};
test_label[3091] = '{-53.8322057263};
test_output[3091] = '{146.37717307};
############ END DEBUG ############*/
test_input[24736:24743] = '{32'h41e6a8b4, 32'h41513dbc, 32'hc20b977a, 32'hc1d8a028, 32'hc28299b4, 32'hc2ac5770, 32'h409dd14b, 32'h4129f5aa};
test_label[3092] = '{32'h409dd14b};
test_output[3092] = '{32'h41bf3462};
/*############ DEBUG ############
test_input[24736:24743] = '{28.8323752282, 13.0775718112, -34.8979258027, -27.0782006705, -65.3002011919, -86.170777997, 4.93179865472, 10.6224769086};
test_label[3092] = '{4.93179865472};
test_output[3092] = '{23.9005767297};
############ END DEBUG ############*/
test_input[24744:24751] = '{32'h42993a08, 32'hc21f8d0f, 32'h41912523, 32'h42997fac, 32'h42c701b4, 32'h427b3a68, 32'h42b767e6, 32'h41b37ec6};
test_label[3093] = '{32'h42993a08};
test_output[3093] = '{32'h41b71f8a};
/*############ DEBUG ############
test_input[24744:24751] = '{76.6133390034, -39.8877532538, 18.1431323913, 76.7493562027, 99.5033301301, 62.8070366491, 91.7029267422, 22.4369006111};
test_label[3093] = '{76.6133390034};
test_output[3093] = '{22.8904006128};
############ END DEBUG ############*/
test_input[24752:24759] = '{32'hc1d78297, 32'h42a5b4b7, 32'hc2792509, 32'h41034583, 32'hc262d6cc, 32'h42b18c2c, 32'hc28c1cde, 32'hc260cee8};
test_label[3094] = '{32'hc28c1cde};
test_output[3094] = '{32'h431ed534};
/*############ DEBUG ############
test_input[24752:24759] = '{-26.938764726, 82.8529577503, -62.2861670995, 8.20447017934, -56.7097626099, 88.7737703174, -70.0563790122, -56.2020567035};
test_label[3094] = '{-70.0563790122};
test_output[3094] = '{158.832828756};
############ END DEBUG ############*/
test_input[24760:24767] = '{32'h41bb99c8, 32'h4094acd7, 32'h422291a7, 32'h426eb420, 32'hc286230b, 32'h428251be, 32'hc299e778, 32'h41f045fb};
test_label[3095] = '{32'h428251be};
test_output[3095] = '{32'h3b87d3f5};
/*############ DEBUG ############
test_input[24760:24767] = '{23.4500880848, 4.64609868436, 40.6422391184, 59.6759045365, -67.0684403819, 65.1596498465, -76.9520859241, 30.0341706497};
test_label[3095] = '{65.1596498465};
test_output[3095] = '{0.00414514051622};
############ END DEBUG ############*/
test_input[24768:24775] = '{32'h42443d07, 32'hc275b642, 32'hc2923d34, 32'hc27e6b8e, 32'h427650f7, 32'hc2267470, 32'h420769c9, 32'hc2a04c8b};
test_label[3096] = '{32'hc2267470};
test_output[3096] = '{32'h42ce62b4};
/*############ DEBUG ############
test_input[24768:24775] = '{49.0595962971, -61.4279849512, -73.1195385058, -63.6050355351, 61.5790660132, -41.613708561, 33.853306726, -80.1494951749};
test_label[3096] = '{-41.613708561};
test_output[3096] = '{103.192778229};
############ END DEBUG ############*/
test_input[24776:24783] = '{32'h425ddfe3, 32'h41d88b2c, 32'h424e2883, 32'hc2575b41, 32'hc218c19c, 32'h422e4d81, 32'hc2c0eb35, 32'h421c5891};
test_label[3097] = '{32'h41d88b2c};
test_output[3097] = '{32'h41e35c7e};
/*############ DEBUG ############
test_input[24776:24783] = '{55.4686400147, 27.0679554363, 51.5395637587, -53.8391159455, -38.1890705728, 43.5756877927, -96.4593869302, 39.0864892611};
test_label[3097] = '{27.0679554363};
test_output[3097] = '{28.4201623901};
############ END DEBUG ############*/
test_input[24784:24791] = '{32'hc2956acb, 32'h42532d7e, 32'hc2a0dc35, 32'h41caf104, 32'h41748137, 32'hc2343256, 32'hc286cbd1, 32'hc2c32d82};
test_label[3098] = '{32'hc286cbd1};
test_output[3098] = '{32'h42f06290};
/*############ DEBUG ############
test_input[24784:24791] = '{-74.7085820846, 52.7944246599, -80.430089355, 25.3676843038, 15.2815461224, -45.0491568241, -67.398080895, -97.5888835906};
test_label[3098] = '{-67.398080895};
test_output[3098] = '{120.192505555};
############ END DEBUG ############*/
test_input[24792:24799] = '{32'hc244f317, 32'hc10df669, 32'h42407343, 32'h42bc4355, 32'h4186472c, 32'hc2842e71, 32'h4216b978, 32'h415dfe3f};
test_label[3099] = '{32'hc10df669};
test_output[3099] = '{32'h42ce0222};
/*############ DEBUG ############
test_input[24792:24799] = '{-49.2373942453, -8.87265864048, 48.1125616732, 94.1315085271, 16.7847513482, -66.0907087088, 37.6811230235, 13.8745715957};
test_label[3099] = '{-8.87265864048};
test_output[3099] = '{103.004167168};
############ END DEBUG ############*/
test_input[24800:24807] = '{32'h42132f6a, 32'h424f1b04, 32'h4223ae6e, 32'hc279ce8b, 32'hc0f48960, 32'hc2526efd, 32'h42bd9581, 32'hc20e944a};
test_label[3100] = '{32'h424f1b04};
test_output[3100] = '{32'h422c0ffe};
/*############ DEBUG ############
test_input[24800:24807] = '{36.7963023576, 51.7763826583, 40.9203419593, -62.4517028924, -7.64176940293, -52.6083872913, 94.7920001033, -35.6448136132};
test_label[3100] = '{51.7763826583};
test_output[3100] = '{43.015617445};
############ END DEBUG ############*/
test_input[24808:24815] = '{32'hc2bae7f6, 32'h4217a4e2, 32'h422f64bb, 32'h41bd512f, 32'h4238c69d, 32'h41ef0cee, 32'hc2831549, 32'hc2a0c756};
test_label[3101] = '{32'h41ef0cee};
test_output[3101] = '{32'h41833c1d};
/*############ DEBUG ############
test_input[24808:24815] = '{-93.4530474235, 37.9110173383, 43.8483680175, 23.6646413669, 46.1939574893, 29.8813125136, -65.5415735722, -80.3893284266};
test_label[3101] = '{29.8813125136};
test_output[3101] = '{16.4043519398};
############ END DEBUG ############*/
test_input[24816:24823] = '{32'h4297cbb7, 32'hc2b4d688, 32'hc25e045c, 32'hc223799c, 32'h423181b2, 32'hc1446150, 32'hc2c66636, 32'h41b3d2fc};
test_label[3102] = '{32'hc1446150};
test_output[3102] = '{32'h42b057e1};
/*############ DEBUG ############
test_input[24816:24823] = '{75.897883249, -90.4190089662, -55.5042584892, -40.8687576831, 44.3766542711, -12.273757921, -99.1996320347, 22.4780200159};
test_label[3102] = '{-12.273757921};
test_output[3102] = '{88.1716411699};
############ END DEBUG ############*/
test_input[24824:24831] = '{32'hc2a2a32b, 32'h41b64c57, 32'h42b2fb92, 32'hc1e2c5a3, 32'h423dcb32, 32'h4237c9d9, 32'hc169674c, 32'hc21bac66};
test_label[3103] = '{32'hc21bac66};
test_output[3103] = '{32'h430068e2};
/*############ DEBUG ############
test_input[24824:24831] = '{-81.3186884211, 22.7872749194, 89.4913464943, -28.3465021897, 47.448434006, 45.9471183601, -14.5877193444, -38.9183570199};
test_label[3103] = '{-38.9183570199};
test_output[3103] = '{128.409703514};
############ END DEBUG ############*/
test_input[24832:24839] = '{32'h419fc451, 32'h425304b2, 32'hc2c24de8, 32'h41bda7b7, 32'h41e20296, 32'h41e4c36e, 32'h428f30b2, 32'h415b454f};
test_label[3104] = '{32'h41bda7b7};
test_output[3104] = '{32'h423f8d88};
/*############ DEBUG ############
test_input[24832:24839] = '{19.9708581328, 52.7545852338, -97.1521642889, 23.7068912704, 28.2512630375, 28.5954253249, 71.5951054652, 13.7044215013};
test_label[3104] = '{23.7068912704};
test_output[3104] = '{47.8882142014};
############ END DEBUG ############*/
test_input[24840:24847] = '{32'hc2b62d1b, 32'h426acf43, 32'h418245b1, 32'hc1866e59, 32'hc2b4112a, 32'hc1aa89cf, 32'h420acdb9, 32'h3e048379};
test_label[3105] = '{32'h3e048379};
test_output[3105] = '{32'h426a4ac0};
/*############ DEBUG ############
test_input[24840:24847] = '{-91.0880987878, 58.7024056679, 16.2840282819, -16.8038815509, -90.0335259802, -21.3172885561, 34.7009013584, 0.12940778181};
test_label[3105] = '{0.12940778181};
test_output[3105] = '{58.5729978861};
############ END DEBUG ############*/
test_input[24848:24855] = '{32'h424c779a, 32'hc2bda7d6, 32'h42b3671d, 32'hc2a4a197, 32'h42c4edb6, 32'hc2702d23, 32'h40a2e526, 32'h40e128ba};
test_label[3106] = '{32'hc2a4a197};
test_output[3106] = '{32'h4334c7b1};
/*############ DEBUG ############
test_input[24848:24855] = '{51.1167969144, -94.8278037015, 89.701389746, -82.3156034684, 98.4642777521, -60.0440774755, 5.09047204292, 7.0362216593};
test_label[3106] = '{-82.3156034684};
test_output[3106] = '{180.78003764};
############ END DEBUG ############*/
test_input[24856:24863] = '{32'h40a37e9c, 32'hc29a5f1a, 32'h4291bcdf, 32'hc242e386, 32'hc2372e0e, 32'hc2807c7f, 32'h41f8a184, 32'h41d86375};
test_label[3107] = '{32'hc29a5f1a};
test_output[3107] = '{32'h43160dfc};
/*############ DEBUG ############
test_input[24856:24863] = '{5.10920546682, -77.1857437728, 72.868889152, -48.7221926885, -45.7949756831, -64.2431595641, 31.0788656027, 27.048562346};
test_label[3107] = '{-77.1857437728};
test_output[3107] = '{150.054632925};
############ END DEBUG ############*/
test_input[24864:24871] = '{32'hc29c1ebe, 32'hc2975ab3, 32'hc21c71e2, 32'h429ced71, 32'hc2c7c2b5, 32'h423b7365, 32'hc20b33e1, 32'h42b9f7c8};
test_label[3108] = '{32'hc21c71e2};
test_output[3108] = '{32'h4304185d};
/*############ DEBUG ############
test_input[24864:24871] = '{-78.060044315, -75.677147545, -39.1112149883, 78.4637520047, -99.8802862495, 46.8626904793, -34.8006627529, 92.9839462605};
test_label[3108] = '{-39.1112149883};
test_output[3108] = '{132.095161743};
############ END DEBUG ############*/
test_input[24872:24879] = '{32'h42782c5f, 32'hc2734790, 32'hc1fa8964, 32'h428ec9c8, 32'h42b43436, 32'hbf42a94c, 32'h42aa5f24, 32'h42ac3b33};
test_label[3109] = '{32'h42b43436};
test_output[3109] = '{32'h3cd16da3};
/*############ DEBUG ############
test_input[24872:24879] = '{62.0433298993, -60.8198849659, -31.3170852735, 71.3941063922, 90.1019740664, -0.760395772569, 85.1858185449, 86.115621146};
test_label[3109] = '{90.1019740664};
test_output[3109] = '{0.0255649743575};
############ END DEBUG ############*/
test_input[24880:24887] = '{32'h41f2ad7f, 32'h42c0dd28, 32'hc26a82af, 32'hc29c416a, 32'h41e410f4, 32'h4284649d, 32'hc233dcc3, 32'h42c465b6};
test_label[3110] = '{32'h41e410f4};
test_output[3110] = '{32'h428bb240};
/*############ DEBUG ############
test_input[24880:24887] = '{30.3347147485, 96.4319423982, -58.6276189414, -78.1277627894, 28.5082774907, 66.1965098525, -44.9655893033, 98.1986558542};
test_label[3110] = '{28.5082774907};
test_output[3110] = '{69.8481456811};
############ END DEBUG ############*/
test_input[24888:24895] = '{32'h42aa66dd, 32'hc2b6ecb4, 32'h42c55758, 32'hc290a33b, 32'h4290468f, 32'h42c1298f, 32'hc2a68e57, 32'hc285c5d7};
test_label[3111] = '{32'h42c55758};
test_output[3111] = '{32'h3deef5ea};
/*############ DEBUG ############
test_input[24888:24895] = '{85.2009068768, -91.4623132659, 98.6705950119, -72.3188088698, 72.1378100772, 96.5811704928, -83.2780060867, -66.8864029847};
test_label[3111] = '{98.6705950119};
test_output[3111] = '{0.116679982223};
############ END DEBUG ############*/
test_input[24896:24903] = '{32'hc287fca0, 32'h41c658f8, 32'h4282537f, 32'hc1bf373e, 32'hc196cb6b, 32'hc1c5cdd3, 32'hc1a6076a, 32'hc25af2ad};
test_label[3112] = '{32'h41c658f8};
test_output[3112] = '{32'h42217a81};
/*############ DEBUG ############
test_input[24896:24903] = '{-67.9934083122, 24.7934418655, 65.1630747887, -23.9019745463, -18.8493261237, -24.7255003121, -20.753620221, -54.7369893921};
test_label[3112] = '{24.7934418655};
test_output[3112] = '{40.3696329232};
############ END DEBUG ############*/
test_input[24904:24911] = '{32'h4278be99, 32'hc25b9fad, 32'hc2a2f7d9, 32'hc2aff62d, 32'h4175b6c5, 32'h422c666a, 32'hc2c57dd0, 32'h42312905};
test_label[3113] = '{32'hc2c57dd0};
test_output[3113] = '{32'h4320ee8e};
/*############ DEBUG ############
test_input[24904:24911] = '{62.1861304251, -54.905933702, -81.4840745287, -87.9808101646, 15.3571212072, 43.1000122594, -98.7457284994, 44.290058334};
test_label[3113] = '{-98.7457284994};
test_output[3113] = '{160.931858947};
############ END DEBUG ############*/
test_input[24912:24919] = '{32'hc1a8808f, 32'hc2079f24, 32'hc21cb412, 32'h42179eed, 32'hc2bd43d9, 32'h42719e8c, 32'h41d0bedd, 32'hc27ee86b};
test_label[3114] = '{32'hc2bd43d9};
test_output[3114] = '{32'h431b098f};
/*############ DEBUG ############
test_input[24912:24919] = '{-21.0627735893, -33.9054112228, -39.1758490706, 37.90520076, -94.6325129907, 60.4048300448, 26.0931940462, -63.7269718945};
test_label[3114] = '{-94.6325129907};
test_output[3114] = '{155.037343036};
############ END DEBUG ############*/
test_input[24920:24927] = '{32'hc13469fa, 32'h42873bcb, 32'hc198581a, 32'h42276cc1, 32'h4259e9b5, 32'hc1280832, 32'hc1d73d4a, 32'hc23acdda};
test_label[3115] = '{32'h4259e9b5};
test_output[3115] = '{32'h41523788};
/*############ DEBUG ############
test_input[24920:24927] = '{-11.2758733269, 67.616786321, -19.0430187695, 41.8562039374, 54.4782303942, -10.502000775, -26.904926017, -46.7010268206};
test_label[3115] = '{54.4782303942};
test_output[3115] = '{13.1385578947};
############ END DEBUG ############*/
test_input[24928:24935] = '{32'hc1c05432, 32'h423c2e50, 32'hc0efaf5e, 32'hc210c721, 32'hc289eeb7, 32'h421b9738, 32'h427089f2, 32'hc2a320e3};
test_label[3116] = '{32'hc2a320e3};
test_output[3116] = '{32'h430db2ee};
/*############ DEBUG ############
test_input[24928:24935] = '{-24.0411106994, 47.045226608, -7.49015705134, -36.1944617406, -68.9662392764, 38.8976737213, 60.1347119573, -81.5642328577};
test_label[3116] = '{-81.5642328577};
test_output[3116] = '{141.698946882};
############ END DEBUG ############*/
test_input[24936:24943] = '{32'hc017cf62, 32'h42765d4d, 32'hc226d39f, 32'hbf9cd9ed, 32'h3f9c5748, 32'hc19b228c, 32'h42c12041, 32'hc1a20e5b};
test_label[3117] = '{32'h42765d4d};
test_output[3117] = '{32'h420be334};
/*############ DEBUG ############
test_input[24936:24943] = '{-2.37203257793, 61.5911137956, -41.7066594904, -1.22540060501, 1.22141362861, -19.3918681573, 96.5629936953, -20.2570100292};
test_label[3117] = '{61.5911137956};
test_output[3117] = '{34.9718798997};
############ END DEBUG ############*/
test_input[24944:24951] = '{32'h4285755b, 32'hc276454c, 32'hc2c2e958, 32'h4292bd41, 32'hc2689b18, 32'hc2116273, 32'h4196cb6e, 32'hc2942ae2};
test_label[3118] = '{32'hc2116273};
test_output[3118] = '{32'h42db6f26};
/*############ DEBUG ############
test_input[24944:24951] = '{66.7292088583, -61.5676736868, -97.4557492322, 73.3696357438, -58.1514570189, -36.3461434556, 18.8493305714, -74.0837528018};
test_label[3118] = '{-36.3461434556};
test_output[3118] = '{109.717084816};
############ END DEBUG ############*/
test_input[24952:24959] = '{32'hc2451156, 32'h42288d44, 32'hc2ae45e2, 32'hc180cd5f, 32'hc23f35a7, 32'hc2b831c4, 32'h41dbf6db, 32'hc24fa034};
test_label[3119] = '{32'hc23f35a7};
test_output[3119] = '{32'h42b3e176};
/*############ DEBUG ############
test_input[24952:24959] = '{-49.266931472, 42.1379545299, -87.1364872749, -16.1002793416, -47.8023947317, -92.0972005311, 27.4955349058, -51.9064475012};
test_label[3119] = '{-47.8023947317};
test_output[3119] = '{89.940349699};
############ END DEBUG ############*/
test_input[24960:24967] = '{32'h42af4e2d, 32'hc298a42d, 32'hc23c874e, 32'hc2b38375, 32'h429077b4, 32'hc247a0e1, 32'hc216a028, 32'h41d7ae83};
test_label[3120] = '{32'h41d7ae83};
test_output[3120] = '{32'h4272c518};
/*############ DEBUG ############
test_input[24960:24967] = '{87.6526841421, -76.3206526465, -47.1321343789, -89.7567533698, 72.2337934601, -49.9071091528, -37.6564025932, 26.9602106887};
test_label[3120] = '{26.9602106887};
test_output[3120] = '{60.6924736547};
############ END DEBUG ############*/
test_input[24968:24975] = '{32'hc22ca1a2, 32'h4277d4f1, 32'hc1ca2faf, 32'hc175e4a1, 32'h42943dcb, 32'hc1332b0e, 32'h41cd08e5, 32'h42485ad1};
test_label[3121] = '{32'h4277d4f1};
test_output[3121] = '{32'h41429a96};
/*############ DEBUG ############
test_input[24968:24975] = '{-43.1578448873, 61.9579507865, -25.2732831472, -15.3683171841, 74.1206863919, -11.1980110699, 25.6293436404, 50.0886877351};
test_label[3121] = '{61.9579507865};
test_output[3121] = '{12.1627408268};
############ END DEBUG ############*/
test_input[24976:24983] = '{32'h42545f39, 32'h42af3a3a, 32'h42b795c5, 32'h40f910c9, 32'h41af463b, 32'h411cab7b, 32'h42579855, 32'hc0a749a0};
test_label[3122] = '{32'h42545f39};
test_output[3122] = '{32'h421adbe3};
/*############ DEBUG ############
test_input[24976:24983] = '{53.0929898655, 87.6137248475, 91.7925223881, 7.78329893674, 21.9092919976, 9.79186519985, 53.8987625021, -5.22773758746};
test_label[3122] = '{53.0929898655};
test_output[3122] = '{38.7147333174};
############ END DEBUG ############*/
test_input[24984:24991] = '{32'h41b1c4bf, 32'hc2aeff44, 32'hc1c698bf, 32'h41b35c90, 32'hc1557a3a, 32'h42c2fdc5, 32'hc26bd84a, 32'h429feb4b};
test_label[3123] = '{32'hc26bd84a};
test_output[3123] = '{32'h431c74f5};
/*############ DEBUG ############
test_input[24984:24991] = '{22.2210678686, -87.4985633553, -24.8245829905, 22.4201964055, -13.3423401641, 97.4956431757, -58.9612198731, 79.9595539104};
test_label[3123] = '{-58.9612198731};
test_output[3123] = '{156.456863073};
############ END DEBUG ############*/
test_input[24992:24999] = '{32'hc2903385, 32'hc2aa0935, 32'hc1b79bf1, 32'h42b25015, 32'hc2c6606c, 32'hc1a70bde, 32'hc1e45f63, 32'hc2036568};
test_label[3124] = '{32'h42b25015};
test_output[3124] = '{32'h80000000};
/*############ DEBUG ############
test_input[24992:24999] = '{-72.1006267458, -85.017985703, -22.9511433748, 89.1564127617, -99.1883274137, -20.8807944617, -28.5465757505, -32.8490277041};
test_label[3124] = '{89.1564127617};
test_output[3124] = '{-0.0};
############ END DEBUG ############*/
test_input[25000:25007] = '{32'h425c4420, 32'h41f672e9, 32'hc268a400, 32'hc2ae4e0e, 32'h4267658b, 32'hc2456c17, 32'hc12a63bf, 32'h429a24be};
test_label[3125] = '{32'hc2456c17};
test_output[3125] = '{32'h42fcdaca};
/*############ DEBUG ############
test_input[25000:25007] = '{55.0665274728, 30.8061089389, -58.1601574012, -87.1524495949, 57.8491627356, -49.3555581861, -10.6493519448, 77.0717642147};
test_label[3125] = '{-49.3555581861};
test_output[3125] = '{126.427322406};
############ END DEBUG ############*/
test_input[25008:25015] = '{32'h42095ba3, 32'hc2a2c727, 32'hc272e79b, 32'hc20b0bd1, 32'hc25e2c5c, 32'hc284e93f, 32'h41229b8e, 32'h42a7e157};
test_label[3126] = '{32'hc272e79b};
test_output[3126] = '{32'h4310aa92};
/*############ DEBUG ############
test_input[25008:25015] = '{34.3394901485, -81.3889675151, -60.7261755303, -34.7615389806, -55.5433214649, -66.4555591568, 10.1629775889, 83.940120284};
test_label[3126] = '{-60.7261755303};
test_output[3126] = '{144.666295814};
############ END DEBUG ############*/
test_input[25016:25023] = '{32'hc25c0ee3, 32'h4213654a, 32'h42b87538, 32'hc239043e, 32'hc2065854, 32'h42bdf158, 32'h4190c3b5, 32'hc1d21406};
test_label[3127] = '{32'hc25c0ee3};
test_output[3127] = '{32'h43160c60};
/*############ DEBUG ############
test_input[25016:25023] = '{-55.0145363321, 36.8489140604, 92.2289460877, -46.2541415178, -33.5862570235, 94.9713738011, 18.0955599781, -26.2597765768};
test_label[3127] = '{-55.0145363321};
test_output[3127] = '{150.048334338};
############ END DEBUG ############*/
test_input[25024:25031] = '{32'h3f8fc031, 32'h418190f0, 32'h4140cba0, 32'h42748334, 32'h4296b316, 32'h41314e2b, 32'hc20b5b6e, 32'hc2afbf27};
test_label[3128] = '{32'h41314e2b};
test_output[3128] = '{32'h42808951};
/*############ DEBUG ############
test_input[25024:25031] = '{1.12305268353, 16.1957708923, 12.049712686, 61.1281288047, 75.3497784232, 11.0815841169, -34.8392868978, -87.873341311};
test_label[3128] = '{11.0815841169};
test_output[3128] = '{64.2681949725};
############ END DEBUG ############*/
test_input[25032:25039] = '{32'h4260ec3b, 32'hc2b20c25, 32'hc2baae7a, 32'h41ea1b71, 32'hc2b7b505, 32'hc298ba15, 32'hc2b5e608, 32'hc1d5f466};
test_label[3129] = '{32'hc1d5f466};
test_output[3129] = '{32'h42a5f337};
/*############ DEBUG ############
test_input[25032:25039] = '{56.2306947404, -89.023718789, -93.340771847, 29.2633988654, -91.8535568667, -76.3634387678, -90.9492818817, -26.7443355257};
test_label[3129] = '{-26.7443355257};
test_output[3129] = '{82.9750302661};
############ END DEBUG ############*/
test_input[25040:25047] = '{32'hc00c2c61, 32'hc1952124, 32'h4201b4f4, 32'h4197c8b3, 32'h429143a1, 32'h42a1064b, 32'h420e3864, 32'hc2058158};
test_label[3130] = '{32'hc00c2c61};
test_output[3130] = '{32'h42a567e0};
/*############ DEBUG ############
test_input[25040:25047] = '{-2.19020871396, -18.6411810342, 32.4267108259, 18.97299779, 72.6320902694, 80.5122934705, 35.5550675339, -33.3763125362};
test_label[3130] = '{-2.19020871396};
test_output[3130] = '{82.7028802692};
############ END DEBUG ############*/
test_input[25048:25055] = '{32'hc1173f4f, 32'hc2255f52, 32'hc29767de, 32'hc2987326, 32'hc29e6439, 32'h42a57046, 32'hc2aa043e, 32'h413abd9c};
test_label[3131] = '{32'hc2987326};
test_output[3131] = '{32'h431ef1b6};
/*############ DEBUG ############
test_input[25048:25055] = '{-9.45295648197, -41.3430846615, -75.7028673439, -76.2249005313, -79.1957478005, 82.7192824422, -85.0082835608, 11.6712912044};
test_label[3131] = '{-76.2249005313};
test_output[3131] = '{158.944182974};
############ END DEBUG ############*/
test_input[25056:25063] = '{32'h42ac69be, 32'hc2b963f6, 32'hc265960f, 32'h42869a19, 32'h41fca6d7, 32'hc2c0fd75, 32'h42810064, 32'hc1d85d18};
test_label[3132] = '{32'hc265960f};
test_output[3132] = '{32'h430f9a63};
/*############ DEBUG ############
test_input[25056:25063] = '{86.2065258285, -92.6952379257, -57.3965414573, 67.3009713546, 31.581464972, -96.4950352891, 64.5007600711, -27.0454550511};
test_label[3132] = '{-57.3965414573};
test_output[3132] = '{143.603067292};
############ END DEBUG ############*/
test_input[25064:25071] = '{32'h428598b8, 32'h42ab2d2f, 32'h41fbc8ed, 32'hc25fa4ae, 32'hc286fa6c, 32'hc0a6de9a, 32'h422a4c1a, 32'h420c88b8};
test_label[3133] = '{32'hc0a6de9a};
test_output[3133] = '{32'h42b59b19};
/*############ DEBUG ############
test_input[25064:25071] = '{66.7982767858, 85.588250029, 31.473107671, -55.910820991, -67.4891066473, -5.21467294871, 42.5743186724, 35.1335139775};
test_label[3133] = '{-5.21467294871};
test_output[3133] = '{90.8029229846};
############ END DEBUG ############*/
test_input[25072:25079] = '{32'h427c47e0, 32'hc003c9cd, 32'h42b43f46, 32'hc28ef466, 32'hc287693a, 32'hc1be924f, 32'hc1576e07, 32'hc26d0647};
test_label[3134] = '{32'hc287693a};
test_output[3134] = '{32'h431dd440};
/*############ DEBUG ############
test_input[25072:25079] = '{63.0701892472, -2.05919200064, 90.1235827174, -71.4773408695, -67.7055219071, -23.821439089, -13.4643625152, -59.2561292776};
test_label[3134] = '{-67.7055219071};
test_output[3134] = '{157.829104624};
############ END DEBUG ############*/
test_input[25080:25087] = '{32'hc1db417f, 32'h42bba11a, 32'hc29eda94, 32'hc1cc0428, 32'h42b353ae, 32'h4242043c, 32'h42b0a969, 32'hc1b7dd29};
test_label[3135] = '{32'h4242043c};
test_output[3135] = '{32'h42355225};
/*############ DEBUG ############
test_input[25080:25087] = '{-27.4069797416, 93.8146523711, -79.4269134485, -25.5020289351, 89.6634397979, 48.5041363668, 88.3308763701, -22.9829892231};
test_label[3135] = '{48.5041363668};
test_output[3135] = '{45.330219537};
############ END DEBUG ############*/
test_input[25088:25095] = '{32'h42b85b62, 32'hc1b5f8a1, 32'h4231ac97, 32'hc2087b9a, 32'h423f55e8, 32'hc22dd5a8, 32'h42b429f5, 32'hc15521f3};
test_label[3136] = '{32'hc22dd5a8};
test_output[3136] = '{32'h4307c0c6};
/*############ DEBUG ############
test_input[25088:25095] = '{92.1784808502, -22.7464011051, 44.4185441342, -34.1207055939, 47.833893781, -43.4586486642, 90.0819455214, -13.3207887805};
test_label[3136] = '{-43.4586486642};
test_output[3136] = '{135.753027606};
############ END DEBUG ############*/
test_input[25096:25103] = '{32'h42b5ae7e, 32'h4134e8d1, 32'hc26b2644, 32'h40610878, 32'hc159e237, 32'h4295f944, 32'hc2a5130b, 32'hc29e1a82};
test_label[3137] = '{32'hc29e1a82};
test_output[3137] = '{32'h4329e480};
/*############ DEBUG ############
test_input[25096:25103] = '{90.840805681, 11.3068396766, -58.7873703678, 3.51614186993, -13.6177280804, 74.9868495121, -82.5371921187, -79.051775602};
test_label[3137] = '{-79.051775602};
test_output[3137] = '{169.892581413};
############ END DEBUG ############*/
test_input[25104:25111] = '{32'h426dd044, 32'h42ab9615, 32'hc23889e3, 32'h42a9e59a, 32'h420accea, 32'hc24d31a3, 32'hc272be95, 32'hc2b7fd51};
test_label[3138] = '{32'h420accea};
test_output[3138] = '{32'h424dcd4a};
/*############ DEBUG ############
test_input[25104:25111] = '{59.453386287, 85.7931305784, -46.1346539351, 84.94844317, 34.7001131699, -51.2984731414, -60.6861163605, -91.9947586823};
test_label[3138] = '{34.7001131699};
test_output[3138] = '{51.4504762038};
############ END DEBUG ############*/
test_input[25112:25119] = '{32'hc28f8253, 32'hc2598b63, 32'hc1d35678, 32'h406eb50a, 32'h423b6fd3, 32'hc2c6662f, 32'hc27ca08d, 32'hc1d4a4dc};
test_label[3139] = '{32'hc27ca08d};
test_output[3139] = '{32'h42dc0830};
/*############ DEBUG ############
test_input[25112:25119] = '{-71.7545401441, -54.3861181998, -26.4172202746, 3.72979976244, 46.8592016373, -99.1995756464, -63.1567880178, -26.5804983836};
test_label[3139] = '{-63.1567880178};
test_output[3139] = '{110.015989655};
############ END DEBUG ############*/
test_input[25120:25127] = '{32'hc1ac6e1f, 32'hbf765bee, 32'h427a975a, 32'hc24665e6, 32'h42336ae7, 32'hc2c5e8ad, 32'h427c8ea6, 32'h428d9697};
test_label[3140] = '{32'h428d9697};
test_output[3140] = '{32'h3a4815fd};
/*############ DEBUG ############
test_input[25120:25127] = '{-21.5537695528, -0.962340241789, 62.6478036512, -49.599510801, 44.8543986494, -98.9544461106, 63.1393049788, 70.7941199163};
test_label[3140] = '{70.7941199163};
test_output[3140] = '{0.000763267104247};
############ END DEBUG ############*/
test_input[25128:25135] = '{32'h41c6a9a2, 32'hc29994f8, 32'h40cf7556, 32'hc25262eb, 32'hc182dd98, 32'h4202d4e7, 32'hc1988075, 32'h42915e08};
test_label[3141] = '{32'h40cf7556};
test_output[3141] = '{32'h428466b3};
/*############ DEBUG ############
test_input[25128:25135] = '{24.8328277247, -76.7909560589, 6.4830730775, -52.5965998008, -16.3581998809, 32.7079141885, -19.0627227558, 72.6836563438};
test_label[3141] = '{6.4830730775};
test_output[3141] = '{66.2005832663};
############ END DEBUG ############*/
test_input[25136:25143] = '{32'h412edbbd, 32'hc0428515, 32'hc28ff4b3, 32'h42ad856f, 32'h4212a491, 32'hc2a5b82e, 32'hbf6c5ee3, 32'hc2195e82};
test_label[3142] = '{32'hc2195e82};
test_output[3142] = '{32'h42fa34b0};
/*############ DEBUG ############
test_input[25136:25143] = '{10.9286471802, -3.03937269124, -71.9779282006, 86.7606152108, 36.6607078412, -82.8597239706, -0.923322860142, -38.3422912443};
test_label[3142] = '{-38.3422912443};
test_output[3142] = '{125.102906455};
############ END DEBUG ############*/
test_input[25144:25151] = '{32'hc2397ab8, 32'h42515b5a, 32'h41f39b0d, 32'hc2172738, 32'h4259367d, 32'h42a9659e, 32'h42b29dac, 32'hc212e95f};
test_label[3143] = '{32'h42b29dac};
test_output[3143] = '{32'h3c225448};
/*############ DEBUG ############
test_input[25144:25151] = '{-46.3698430819, 52.3392122409, 30.4507075214, -37.7883009043, 54.3032127571, 84.6984746731, 89.3079506966, -36.7278995682};
test_label[3143] = '{89.3079506966};
test_output[3143] = '{0.00990778954552};
############ END DEBUG ############*/
test_input[25152:25159] = '{32'h41c63be8, 32'h41004329, 32'h4165acf7, 32'hc1a0e2f3, 32'h4280a2ba, 32'hc28044cf, 32'hc0f4ba6b, 32'hc29b26a6};
test_label[3144] = '{32'hc1a0e2f3};
test_output[3144] = '{32'h42a8db77};
/*############ DEBUG ############
test_input[25152:25159] = '{24.7792510261, 8.01639626919, 14.3547274344, -20.1108149899, 64.317823783, -64.1343915345, -7.64775604258, -77.5754826223};
test_label[3144] = '{-20.1108149899};
test_output[3144] = '{84.428638773};
############ END DEBUG ############*/
test_input[25160:25167] = '{32'hc29c22ca, 32'hc28b3aec, 32'h428f25e2, 32'h417867b0, 32'hc23edf7e, 32'hc25338c1, 32'hc1cf02c2, 32'h42b6b548};
test_label[3145] = '{32'h428f25e2};
test_output[3145] = '{32'h419e3d98};
/*############ DEBUG ############
test_input[25160:25167] = '{-78.0679498343, -69.6150799882, 71.5739930688, 15.5253141506, -47.7182549367, -52.8054249901, -25.8763461108, 91.3540673638};
test_label[3145] = '{71.5739930688};
test_output[3145] = '{19.7800742976};
############ END DEBUG ############*/
test_input[25168:25175] = '{32'h42c32543, 32'hc10e41a8, 32'h429a4511, 32'hc2c7a265, 32'hc228be4a, 32'hc1825e4d, 32'hc13bde36, 32'h427cdc69};
test_label[3146] = '{32'hc13bde36};
test_output[3146] = '{32'h42daa109};
/*############ DEBUG ############
test_input[25168:25175] = '{97.5727732465, -8.89102967711, 77.1348939891, -99.8171781273, -42.1858299835, -16.2960446629, -11.7417506247, 63.215245495};
test_label[3146] = '{-11.7417506247};
test_output[3146] = '{109.314523873};
############ END DEBUG ############*/
test_input[25176:25183] = '{32'h4238ac85, 32'hc2399b6a, 32'hc2bcb191, 32'h425d960a, 32'hc2a0b27c, 32'h417b7d5e, 32'hc22de937, 32'h4187e13b};
test_label[3147] = '{32'hc22de937};
test_output[3147] = '{32'h42c5bfae};
/*############ DEBUG ############
test_input[25176:25183] = '{46.1684770062, -46.4017698315, -94.3468091451, 55.3965243918, -80.348599228, 15.7181074084, -43.4777488044, 16.9849764545};
test_label[3147] = '{-43.4777488044};
test_output[3147] = '{98.8743714362};
############ END DEBUG ############*/
test_input[25184:25191] = '{32'hc2a18c90, 32'h42a8cf31, 32'hc2a62307, 32'hc299ef22, 32'hc29830a2, 32'hc2826e64, 32'h423a72d8, 32'hc26f56bd};
test_label[3148] = '{32'h423a72d8};
test_output[3148] = '{32'h42172b8a};
/*############ DEBUG ############
test_input[25184:25191] = '{-80.7745398516, 84.4046715369, -83.0684098193, -76.9670554899, -76.0949829899, -65.2156070072, 46.6121538391, -59.8347051335};
test_label[3148] = '{46.6121538391};
test_output[3148] = '{37.7925176978};
############ END DEBUG ############*/
test_input[25192:25199] = '{32'h42b4ccf5, 32'h4267556a, 32'hc2055eba, 32'hc1f16cca, 32'h41e4b9c5, 32'hc273e9c5, 32'h428bdefe, 32'h422331a4};
test_label[3149] = '{32'hc273e9c5};
test_output[3149] = '{32'h431760ec};
/*############ DEBUG ############
test_input[25192:25199] = '{90.4003071806, 57.8334133237, -33.3425055746, -30.1781188237, 28.590708635, -60.9782902017, 69.93553463, 40.7984754801};
test_label[3149] = '{-60.9782902017};
test_output[3149] = '{151.378597384};
############ END DEBUG ############*/
test_input[25200:25207] = '{32'h42b90ea7, 32'h42619b80, 32'hc26307d0, 32'h42a233fb, 32'hc211344f, 32'hc22a8621, 32'hc21891a2, 32'hc23f925c};
test_label[3150] = '{32'hc22a8621};
test_output[3150] = '{32'h430728dc};
/*############ DEBUG ############
test_input[25200:25207] = '{92.5286195945, 56.4018557729, -56.7576276505, 81.1015217778, -36.3010829409, -42.630983458, -38.142218043, -47.8929271935};
test_label[3150] = '{-42.630983458};
test_output[3150] = '{135.159613949};
############ END DEBUG ############*/
test_input[25208:25215] = '{32'hc2222c07, 32'hc1e90b6f, 32'h42aa6fe5, 32'h40622d37, 32'hc2c5565f, 32'h4138c5f0, 32'hc2b244ba, 32'hc291e34c};
test_label[3151] = '{32'hc2222c07};
test_output[3151] = '{32'h42fb85e8};
/*############ DEBUG ############
test_input[25208:25215] = '{-40.5429950256, -29.1305833896, 85.2185407238, 3.53400961243, -98.6686899624, 11.5483243175, -89.1342322376, -72.9439423742};
test_label[3151] = '{-40.5429950256};
test_output[3151] = '{125.761535749};
############ END DEBUG ############*/
test_input[25216:25223] = '{32'hc2801c97, 32'h42778b65, 32'h42abb8a8, 32'h4202a201, 32'h4246b334, 32'hc2c183fe, 32'hc291c7bf, 32'hc290d5b9};
test_label[3152] = '{32'hc290d5b9};
test_output[3152] = '{32'h431e4730};
/*############ DEBUG ############
test_input[25216:25223] = '{-64.0558384714, 61.8861279657, 85.8606545887, 32.6582073247, 49.6750048988, -96.757794253, -72.8901290663, -72.4174234358};
test_label[3152] = '{-72.4174234358};
test_output[3152] = '{158.278078024};
############ END DEBUG ############*/
test_input[25224:25231] = '{32'hc266b595, 32'h41223686, 32'hc25c6e0f, 32'hc2bac2e9, 32'hc2749241, 32'hc24110bf, 32'hc2bfa383, 32'h420e4eeb};
test_label[3153] = '{32'hc25c6e0f};
test_output[3153] = '{32'h42b55e7d};
/*############ DEBUG ############
test_input[25224:25231] = '{-57.6773254307, 10.1383110344, -55.1074776522, -93.3806872038, -61.1428244611, -48.2663546681, -95.8193560729, 35.5770679893};
test_label[3153] = '{-55.1074776522};
test_output[3153] = '{90.6845456415};
############ END DEBUG ############*/
test_input[25232:25239] = '{32'h42880a45, 32'h4228b213, 32'h42909f24, 32'hc0826ccd, 32'hc2610dc8, 32'hc1ba1ce6, 32'h426f1d88, 32'hc2552755};
test_label[3154] = '{32'hc2610dc8};
test_output[3154] = '{32'h43009680};
/*############ DEBUG ############
test_input[25232:25239] = '{68.0200581349, 42.173899637, 72.3108241455, -4.0757815536, -56.2634577131, -23.2641112357, 59.7788373538, -53.288409126};
test_label[3154] = '{-56.2634577131};
test_output[3154] = '{128.587886929};
############ END DEBUG ############*/
test_input[25240:25247] = '{32'h4137d165, 32'hc1acf245, 32'h42ba1ef4, 32'hc22f8260, 32'h429d8241, 32'h429ba4bd, 32'hc184297c, 32'hbf3386c9};
test_label[3155] = '{32'hc184297c};
test_output[3155] = '{32'h42db2953};
/*############ DEBUG ############
test_input[25240:25247] = '{11.4886217894, -21.6182961362, 93.0604528763, -43.87731934, 78.7544045815, 77.8217565815, -16.5202569591, -0.701275425056};
test_label[3155] = '{-16.5202569591};
test_output[3155] = '{109.580710689};
############ END DEBUG ############*/
test_input[25248:25255] = '{32'hc25a9f9c, 32'h420e0232, 32'hc28ab59b, 32'hc1e6a1a4, 32'h42035881, 32'h429b5323, 32'hc2944671, 32'hc2113835};
test_label[3156] = '{32'hc2944671};
test_output[3156] = '{32'h4317ccca};
/*############ DEBUG ############
test_input[25248:25255] = '{-54.6558689064, 35.5021438022, -69.3546971348, -28.8289256976, 32.8364290567, 77.6623751012, -74.1375790638, -36.3048884775};
test_label[3156] = '{-74.1375790638};
test_output[3156] = '{151.799954165};
############ END DEBUG ############*/
test_input[25256:25263] = '{32'h3f037eba, 32'hc0000d4e, 32'hc283b6bf, 32'hc1e2f285, 32'hc28c581b, 32'hc0ea251f, 32'hc2867be6, 32'hc288f990};
test_label[3157] = '{32'hc2867be6};
test_output[3157] = '{32'h4287aae9};
/*############ DEBUG ############
test_input[25256:25263] = '{0.51365244497, -2.00081193873, -65.8569254523, -28.3684168397, -70.1720776556, -7.31703156515, -67.2419906736, -68.4874295851};
test_label[3157] = '{-67.2419906736};
test_output[3157] = '{67.8338104586};
############ END DEBUG ############*/
test_input[25264:25271] = '{32'hc2a2b589, 32'hc29082c0, 32'hc10d9d7b, 32'h401cd7fd, 32'h409836dc, 32'h424a00bd, 32'h42b49d05, 32'h429f8e01};
test_label[3158] = '{32'h429f8e01};
test_output[3158] = '{32'h4128783c};
/*############ DEBUG ############
test_input[25264:25271] = '{-81.3545625233, -72.2553747648, -8.85094700699, 2.45068288623, 4.75669657981, 50.5007217405, 90.3066756977, 79.7773482615};
test_label[3158] = '{79.7773482615};
test_output[3158] = '{10.5293541765};
############ END DEBUG ############*/
test_input[25272:25279] = '{32'h420e52ee, 32'hc2a634d7, 32'hc296ef9a, 32'hc1a1d290, 32'h4247e90a, 32'hc20e32da, 32'hc264cc0e, 32'hc12ef7af};
test_label[3159] = '{32'hc296ef9a};
test_output[3159] = '{32'h42fae41e};
/*############ DEBUG ############
test_input[25272:25279] = '{35.5809865254, -83.1032032054, -75.4679682129, -20.2278144287, 49.9775758374, -35.5496603574, -57.1992737417, -10.9354697769};
test_label[3159] = '{-75.4679682129};
test_output[3159] = '{125.44554461};
############ END DEBUG ############*/
test_input[25280:25287] = '{32'hc28475d4, 32'h41942d97, 32'h41a5f8ab, 32'hc26904d8, 32'hc2a22f8e, 32'h40bfd5ac, 32'hc248fbd4, 32'hc190f5c4};
test_label[3160] = '{32'h40bfd5ac};
test_output[3160] = '{32'h416dab29};
/*############ DEBUG ############
test_input[25280:25287] = '{-66.230135554, 18.5222603575, 20.7464206909, -58.2547319977, -81.0928781523, 5.99483286191, -50.2459258015, -18.1200020545};
test_label[3160] = '{5.99483286191};
test_output[3160] = '{14.8542875384};
############ END DEBUG ############*/
test_input[25288:25295] = '{32'hc28e6ee8, 32'hc2c43340, 32'hc1bf7720, 32'hc1a9c902, 32'h424cc7ba, 32'hc2a4118e, 32'h4295f49e, 32'hc20b18ab};
test_label[3161] = '{32'hc2c43340};
test_output[3161] = '{32'h432d13ef};
/*############ DEBUG ############
test_input[25288:25295] = '{-71.2166141397, -98.1000960988, -23.93316658, -21.2231480582, 51.1950457441, -82.0342875414, 74.9777714627, -34.7740916424};
test_label[3161] = '{-98.1000960988};
test_output[3161] = '{173.077867562};
############ END DEBUG ############*/
test_input[25296:25303] = '{32'h42a83bb0, 32'h40a8ce32, 32'hc213e499, 32'hc1dbbae1, 32'hc2be2283, 32'h429ba359, 32'h405ebb9c, 32'hc2957da7};
test_label[3162] = '{32'h42a83bb0};
test_output[3162] = '{32'h3af10eea};
/*############ DEBUG ############
test_input[25296:25303] = '{84.1165790825, 5.27517028798, -36.9732384858, -27.4662502325, -95.0674048665, 77.8190353508, 3.48020070538, -74.7454139602};
test_label[3162] = '{84.1165790825};
test_output[3162] = '{0.00183912854404};
############ END DEBUG ############*/
test_input[25304:25311] = '{32'hc27d53e0, 32'h42885cdd, 32'h41f28def, 32'hc27a3a73, 32'hc1832ec5, 32'hc2891dd7, 32'hc2abcfbb, 32'h4294d4c7};
test_label[3163] = '{32'hc27a3a73};
test_output[3163] = '{32'h4308f981};
/*############ DEBUG ############
test_input[25304:25311] = '{-63.3319096989, 68.1813748826, 30.3193030863, -62.5570789221, -16.3978370932, -68.5582837302, -85.9057247609, 74.415581613};
test_label[3163] = '{-62.5570789221};
test_output[3163] = '{136.974619799};
############ END DEBUG ############*/
test_input[25312:25319] = '{32'h4185b4d4, 32'h413154c2, 32'h41a5e0d1, 32'h42466038, 32'hc27a308a, 32'hc1f4d651, 32'hc2b29e30, 32'h42a7701f};
test_label[3164] = '{32'hc27a308a};
test_output[3164] = '{32'h43124432};
/*############ DEBUG ############
test_input[25312:25319] = '{16.7132944258, 11.0831928519, 20.7347733362, 49.5939636442, -62.5474006286, -30.6046474539, -89.3089567957, 83.7189848343};
test_label[3164] = '{-62.5474006286};
test_output[3164] = '{146.266385463};
############ END DEBUG ############*/
test_input[25320:25327] = '{32'hc1c90a3e, 32'h418204c2, 32'h427058dd, 32'h425b9132, 32'hc2547d19, 32'hc2c7b75c, 32'h42398e85, 32'h4259f10e};
test_label[3165] = '{32'hc1c90a3e};
test_output[3165] = '{32'h42aa73b3};
/*############ DEBUG ############
test_input[25320:25327] = '{-25.1300017253, 16.252323448, 60.0867792777, 54.8917922797, -53.1221660717, -99.8581274717, 46.3891773382, 54.4854055128};
test_label[3165] = '{-25.1300017253};
test_output[3165] = '{85.2259767926};
############ END DEBUG ############*/
test_input[25328:25335] = '{32'h42acd732, 32'h42aa0e95, 32'hc290ea14, 32'h40df9dea, 32'hc2052054, 32'hc2930c51, 32'hc11d2dde, 32'hbf3034a5};
test_label[3166] = '{32'hc2930c51};
test_output[3166] = '{32'h43202a99};
/*############ DEBUG ############
test_input[25328:25335] = '{86.4203057581, 85.0284776768, -72.4571807953, 6.98802667724, -33.2815710864, -73.5240545422, -9.8236976979, -0.688303314503};
test_label[3166] = '{-73.5240545422};
test_output[3166] = '{160.166399555};
############ END DEBUG ############*/
test_input[25336:25343] = '{32'hc281327a, 32'hc1b2ee9a, 32'hc28915d6, 32'hc0c8f0b9, 32'h420e03e0, 32'hc207a24e, 32'h4295838e, 32'hc2bcc9f6};
test_label[3167] = '{32'hc2bcc9f6};
test_output[3167] = '{32'h432926c2};
/*############ DEBUG ############
test_input[25336:25343] = '{-64.5985867112, -22.3665048109, -68.5426452253, -6.27938506561, 35.5037823747, -33.9084999959, 74.7569450337, -94.3944518183};
test_label[3167] = '{-94.3944518183};
test_output[3167] = '{169.151396852};
############ END DEBUG ############*/
test_input[25344:25351] = '{32'h42aaacaf, 32'hc1d80c48, 32'hc22ef48d, 32'hc2226af6, 32'hc221ff12, 32'h41d2cb3a, 32'h427c6116, 32'hc22e4b3a};
test_label[3168] = '{32'hc1d80c48};
test_output[3168] = '{32'h42e0afc1};
/*############ DEBUG ############
test_input[25344:25351] = '{85.3372717636, -27.0059968205, -43.738819568, -40.6044531237, -40.4990904933, 26.3492314223, 63.0948115787, -43.5734631243};
test_label[3168] = '{-27.0059968205};
test_output[3168] = '{112.343268584};
############ END DEBUG ############*/
test_input[25352:25359] = '{32'hc2483358, 32'hc2a0051a, 32'h42752b92, 32'hc2b48ab6, 32'h42a86e79, 32'h429f9ff2, 32'h41ad0800, 32'hc2b3b583};
test_label[3169] = '{32'hc2b3b583};
test_output[3169] = '{32'h432e151b};
/*############ DEBUG ############
test_input[25352:25359] = '{-50.0501415425, -80.0099648229, 61.292548844, -90.2709235639, 84.21576663, 79.812393314, 21.6289058427, -89.8545123871};
test_label[3169] = '{-89.8545123871};
test_output[3169] = '{174.082440757};
############ END DEBUG ############*/
test_input[25360:25367] = '{32'hc1db861e, 32'hc1f913dc, 32'hc23dffe4, 32'hc266b28d, 32'hc26dfe4a, 32'h41d7760f, 32'h419d5e05, 32'h42b65e72};
test_label[3170] = '{32'h41d7760f};
test_output[3170] = '{32'h428080ee};
/*############ DEBUG ############
test_input[25360:25367] = '{-27.4404873856, -31.1346974783, -47.4998930618, -57.6743667629, -59.4983284908, 26.9326453808, 19.6709085003, 91.1844609507};
test_label[3170] = '{26.9326453808};
test_output[3170] = '{64.2518155699};
############ END DEBUG ############*/
test_input[25368:25375] = '{32'h41b1a3b6, 32'hc2a744f0, 32'hc18b635c, 32'h422c9003, 32'hc1054bf2, 32'h42ad03ae, 32'hc2b6d500, 32'h4285663f};
test_label[3171] = '{32'h4285663f};
test_output[3171] = '{32'h419e75bc};
/*############ DEBUG ############
test_input[25368:25375] = '{22.2049361137, -83.6346452626, -17.4235146987, 43.1406378348, -8.33104088308, 86.5071884428, -91.4160175148, 66.6997014531};
test_label[3171] = '{66.6997014531};
test_output[3171] = '{19.8074869922};
############ END DEBUG ############*/
test_input[25376:25383] = '{32'h42a35408, 32'hc22472c1, 32'hc27e3606, 32'hc296f214, 32'h421a8eb8, 32'h42547cc1, 32'hc1b96ca8, 32'hc217923c};
test_label[3172] = '{32'hc27e3606};
test_output[3172] = '{32'h43113786};
/*############ DEBUG ############
test_input[25376:25383] = '{81.6641250489, -41.1120642933, -63.5527588608, -75.4728078383, 38.6393742073, 53.1218290698, -23.1780541988, -37.8928064094};
test_label[3172] = '{-63.5527588608};
test_output[3172] = '{145.21688391};
############ END DEBUG ############*/
test_input[25384:25391] = '{32'hc21e9a03, 32'hc1defc98, 32'h42aeca50, 32'h4238dcb6, 32'hc29ab79d, 32'h425ea785, 32'hc1fc9cd8, 32'h42994154};
test_label[3173] = '{32'hc1fc9cd8};
test_output[3173] = '{32'h42edf188};
/*############ DEBUG ############
test_input[25384:25391] = '{-39.6504031842, -27.8733370692, 87.3951385222, 46.215537955, -77.3586234425, 55.6635935995, -31.5765839332, 76.6275927721};
test_label[3173] = '{-31.5765839332};
test_output[3173] = '{118.971743528};
############ END DEBUG ############*/
test_input[25392:25399] = '{32'h4263e230, 32'hc2b0e83b, 32'hc2804ae8, 32'hc2219653, 32'hc27d69b0, 32'h427189f4, 32'h422e0b20, 32'h4214d9a6};
test_label[3174] = '{32'hc2804ae8};
test_output[3174] = '{32'h42f92077};
/*############ DEBUG ############
test_input[25392:25399] = '{56.9708851154, -88.4535729136, -64.1463036006, -40.3968013343, -63.3532086256, 60.3847205516, 43.5108651314, 37.2125464011};
test_label[3174] = '{-64.1463036006};
test_output[3174] = '{124.563408825};
############ END DEBUG ############*/
test_input[25400:25407] = '{32'hc10f7c2c, 32'hc21feebc, 32'h428e3b46, 32'hc27e9da5, 32'h42838682, 32'hc2805793, 32'h42421a15, 32'h424f5d58};
test_label[3175] = '{32'h424f5d58};
test_output[3175] = '{32'h419a3c14};
/*############ DEBUG ############
test_input[25400:25407] = '{-8.96781549521, -39.9831407223, 71.1157703018, -63.6539509138, 65.7627117436, -64.1710421251, 48.5254719407, 51.841157354};
test_label[3175] = '{51.841157354};
test_output[3175] = '{19.2793354344};
############ END DEBUG ############*/
test_input[25408:25415] = '{32'hc29c6c60, 32'h42187487, 32'h42923c37, 32'h42c41a83, 32'h409af950, 32'h42a99ed0, 32'h422012fa, 32'hc299875f};
test_label[3176] = '{32'h409af950};
test_output[3176] = '{32'h42ba6aee};
/*############ DEBUG ############
test_input[25408:25415] = '{-78.2116680186, 38.1137961632, 73.1176073791, 98.0517826031, 4.84293364359, 84.8101806883, 40.0185328904, -76.76439382};
test_label[3176] = '{4.84293364359};
test_output[3176] = '{93.2088507347};
############ END DEBUG ############*/
test_input[25416:25423] = '{32'hc1f05f4e, 32'hc1bf415c, 32'hc242ce9c, 32'h41e87980, 32'hc0e11ebd, 32'hc222a9a2, 32'h4019b33c, 32'h4286e928};
test_label[3177] = '{32'hc222a9a2};
test_output[3177] = '{32'h42d83df9};
/*############ DEBUG ############
test_input[25416:25423] = '{-30.0465353436, -23.9069133514, -48.7017688169, 29.0593261275, -7.03500214928, -40.6656558064, 2.40156463287, 67.4553807626};
test_label[3177] = '{-40.6656558064};
test_output[3177] = '{108.121036569};
############ END DEBUG ############*/
test_input[25424:25431] = '{32'h41c4b13a, 32'hc2865fa1, 32'h42194b96, 32'hc13c9d0c, 32'hc1e33801, 32'hc2832808, 32'h40daa71c, 32'h420b19f4};
test_label[3178] = '{32'hc2865fa1};
test_output[3178] = '{32'h42d313f2};
/*############ DEBUG ############
test_input[25424:25431] = '{24.5865368486, -67.1867763529, 38.3238130082, -11.7883416578, -28.4023457385, -65.5781851895, 6.83289911423, 34.7753437373};
test_label[3178] = '{-67.1867763529};
test_output[3178] = '{105.538953007};
############ END DEBUG ############*/
test_input[25432:25439] = '{32'h3fc54609, 32'hc18fb42c, 32'hc1087134, 32'h42ae4bfd, 32'h429dc6f1, 32'h4220a644, 32'hc1b8d0e4, 32'hc2aed37e};
test_label[3179] = '{32'hc1087134};
test_output[3179] = '{32'h42bf5a45};
/*############ DEBUG ############
test_input[25432:25439] = '{1.54119981085, -17.9629740568, -8.52763720769, 87.1484146267, 78.8885598114, 40.1623701715, -23.1019978551, -87.4130689267};
test_label[3179] = '{-8.52763720769};
test_output[3179] = '{95.6763104975};
############ END DEBUG ############*/
test_input[25440:25447] = '{32'hc2836f27, 32'h42a1815d, 32'hc25caf2e, 32'h4256c7c9, 32'h42ae870f, 32'hc147a658, 32'h42b205b0, 32'h42a96738};
test_label[3180] = '{32'h42a96738};
test_output[3180] = '{32'h408f6a54};
/*############ DEBUG ############
test_input[25440:25447] = '{-65.717094725, 80.7526612664, -55.1710743388, 53.6951042221, 87.2637851042, -12.4781110978, 89.0111050059, 84.7015955565};
test_label[3180] = '{84.7015955565};
test_output[3180] = '{4.48172974506};
############ END DEBUG ############*/
test_input[25448:25455] = '{32'h41a7a36a, 32'hc2337dc6, 32'h420fc448, 32'h42b5007b, 32'h416855f5, 32'h4282f4ff, 32'hc1714252, 32'h42953962};
test_label[3181] = '{32'h41a7a36a};
test_output[3181] = '{32'h428b17a1};
/*############ DEBUG ############
test_input[25448:25455] = '{20.9547914179, -44.8728243432, 35.9416801807, 90.5009400093, 14.5209855623, 65.4785043071, -15.0786913455, 74.6120768148};
test_label[3181] = '{20.9547914179};
test_output[3181] = '{69.5461487172};
############ END DEBUG ############*/
test_input[25456:25463] = '{32'h42b4d97b, 32'hc22ed6d3, 32'hc2354d2d, 32'h42bc98d7, 32'hc14b4a92, 32'hc2117519, 32'hc24aaf81, 32'hc046622a};
test_label[3182] = '{32'h42b4d97b};
test_output[3182] = '{32'h40793c7d};
/*############ DEBUG ############
test_input[25456:25463] = '{90.424766752, -43.7097911532, -45.3253671113, 94.2985164109, -12.7057056265, -36.3643514305, -50.6713915704, -3.09974157481};
test_label[3182] = '{90.424766752};
test_output[3182] = '{3.89431699774};
############ END DEBUG ############*/
test_input[25464:25471] = '{32'hc29408c8, 32'hc0ea4c0c, 32'h3f8b5287, 32'h42be157a, 32'h41e14de3, 32'h41409d98, 32'hc2592309, 32'h42800777};
test_label[3183] = '{32'hc29408c8};
test_output[3183] = '{32'h43290f21};
/*############ DEBUG ############
test_input[25464:25471] = '{-74.0171502072, -7.32178286294, 1.08845598359, 95.0419468078, 28.1630310122, 12.0384747524, -54.2842135346, 64.0145819284};
test_label[3183] = '{-74.0171502072};
test_output[3183] = '{169.059097015};
############ END DEBUG ############*/
test_input[25472:25479] = '{32'h42a45631, 32'hc1406066, 32'hc220bd8e, 32'hc1a08871, 32'h42ad22bb, 32'h42bc1c0c, 32'hc1383590, 32'h42a4600f};
test_label[3184] = '{32'h42bc1c0c};
test_output[3184] = '{32'h3a167e7b};
/*############ DEBUG ############
test_input[25472:25479] = '{82.1683389824, -12.0235347867, -40.1851101982, -20.0666211573, 86.5678345272, 94.0547765795, -11.5130768067, 82.18761399};
test_label[3184] = '{94.0547765795};
test_output[3184] = '{0.000574089267194};
############ END DEBUG ############*/
test_input[25480:25487] = '{32'h42734a79, 32'hc175befb, 32'hc1d3d406, 32'h418f2e3e, 32'hc164a02f, 32'h42c778e9, 32'hc27212cd, 32'h40d77fb9};
test_label[3185] = '{32'hc1d3d406};
test_output[3185] = '{32'h42fc6deb};
/*############ DEBUG ############
test_input[25480:25487] = '{60.8227262303, -15.3591262519, -26.4785272813, 17.8975797116, -14.289107455, 99.7361532225, -60.5183617945, 6.73434128447};
test_label[3185] = '{-26.4785272813};
test_output[3185] = '{126.214680504};
############ END DEBUG ############*/
test_input[25488:25495] = '{32'h4027c976, 32'h4201f340, 32'h4285d683, 32'hc0932d4b, 32'hc090fdcf, 32'hc1faeae7, 32'hc2a3a910, 32'h42bb84a3};
test_label[3186] = '{32'hc090fdcf};
test_output[3186] = '{32'h42c49480};
/*############ DEBUG ############
test_input[25488:25495] = '{2.62167116288, 32.487547175, 66.9189670918, -4.59927887733, -4.53098269136, -31.364697581, -81.8302015376, 93.7590557935};
test_label[3186] = '{-4.53098269136};
test_output[3186] = '{98.2900384848};
############ END DEBUG ############*/
test_input[25496:25503] = '{32'hc24dafb6, 32'hbfeb6af9, 32'h42649d2f, 32'h41169c69, 32'h41e22984, 32'hc211db25, 32'hc1f65507, 32'h429cbc4d};
test_label[3187] = '{32'hc1f65507};
test_output[3187] = '{32'h42da518e};
/*############ DEBUG ############
test_input[25496:25503] = '{-51.4215924595, -1.83920202411, 57.1534988754, 9.4131864614, 28.2702712807, -36.4640084174, -30.791517204, 78.3677719421};
test_label[3187] = '{-30.791517204};
test_output[3187] = '{109.159289147};
############ END DEBUG ############*/
test_input[25504:25511] = '{32'h42061e55, 32'hc241f51b, 32'h42b98d28, 32'hc2470c1c, 32'hc2849583, 32'h420fcfdc, 32'hc2524419, 32'h418a9d8a};
test_label[3188] = '{32'hc2470c1c};
test_output[3188] = '{32'h430e899b};
/*############ DEBUG ############
test_input[25504:25511] = '{33.5296228672, -48.4893624761, 92.7756976881, -49.7618254399, -66.2920130947, 35.9529876749, -52.5665010594, 17.3269233626};
test_label[3188] = '{-49.7618254399};
test_output[3188] = '{142.537523128};
############ END DEBUG ############*/
test_input[25512:25519] = '{32'hc28991e8, 32'hc2bcf89e, 32'h40c82903, 32'hc2126564, 32'h42c5cd91, 32'hc1b158cf, 32'hc21ebd6f, 32'h41563229};
test_label[3189] = '{32'h41563229};
test_output[3189] = '{32'h42ab074c};
/*############ DEBUG ############
test_input[25512:25519] = '{-68.7849729808, -94.4855832247, 6.25500628882, -36.5990127758, 98.9014965011, -22.1683634528, -39.6849927059, 13.3872463363};
test_label[3189] = '{13.3872463363};
test_output[3189] = '{85.5142501648};
############ END DEBUG ############*/
test_input[25520:25527] = '{32'h42c37a01, 32'hc14d4b6f, 32'h42c103fb, 32'hc2c29354, 32'h417877ac, 32'h40ef6fa6, 32'hc24b21b2, 32'h428847cd};
test_label[3190] = '{32'h428847cd};
test_output[3190] = '{32'h41eed5b7};
/*############ DEBUG ############
test_input[25520:25527] = '{97.7382886893, -12.8309167209, 96.5077705834, -97.2877524316, 15.5292168344, 7.48237890905, -50.7829041382, 68.1402372294};
test_label[3190] = '{68.1402372294};
test_output[3190] = '{29.8543521305};
############ END DEBUG ############*/
test_input[25528:25535] = '{32'hc2a3871c, 32'h4176d21f, 32'h427c11f7, 32'h42743070, 32'h4290a254, 32'hc2a25333, 32'h415c81b6, 32'hc1e80cc0};
test_label[3191] = '{32'h415c81b6};
test_output[3191] = '{32'h426a2456};
/*############ DEBUG ############
test_input[25528:25535] = '{-81.7638842075, 15.4262986951, 63.0175449306, 61.0473008447, 72.317047534, -81.1625017249, 13.7816673751, -29.0062257032};
test_label[3191] = '{13.7816673751};
test_output[3191] = '{58.5354843761};
############ END DEBUG ############*/
test_input[25536:25543] = '{32'hc26b8ef4, 32'hc22b2454, 32'h426fece6, 32'h41361db8, 32'hc25371a2, 32'hc20ce396, 32'h41295d5c, 32'h42a26da1};
test_label[3192] = '{32'hc20ce396};
test_output[3192] = '{32'h42e8df6c};
/*############ DEBUG ############
test_input[25536:25543] = '{-58.8896028412, -42.7854771187, 59.9813479241, 11.3822553878, -52.8609686719, -35.2222505941, 10.5852931244, 81.2141218746};
test_label[3192] = '{-35.2222505941};
test_output[3192] = '{116.436372469};
############ END DEBUG ############*/
test_input[25544:25551] = '{32'hc2256cf2, 32'h41b5f5c2, 32'h428ef615, 32'hc2106951, 32'hc1e2fe10, 32'hc28e6e50, 32'h4252e09c, 32'hc16f8cf5};
test_label[3193] = '{32'h428ef615};
test_output[3193] = '{32'h31f46a35};
/*############ DEBUG ############
test_input[25544:25551] = '{-41.3563914822, 22.7449993127, 71.480629812, -36.1028476138, -28.3740533369, -71.2154543596, 52.7193455524, -14.9719134342};
test_label[3193] = '{71.480629812};
test_output[3193] = '{7.11340888725e-09};
############ END DEBUG ############*/
test_input[25552:25559] = '{32'hc21c18dd, 32'h42ae7795, 32'hc206f57a, 32'h3ed3908d, 32'hc2c12062, 32'h4285d76b, 32'h42ab624d, 32'hc27c161b};
test_label[3194] = '{32'h42ae7795};
test_output[3194] = '{32'h3e469ce3};
/*############ DEBUG ############
test_input[25552:25559] = '{-39.0242815678, 87.2335594005, -33.7397230324, 0.413212213032, -96.5632463395, 66.9207386574, 85.6919908881, -63.021587621};
test_label[3194] = '{87.2335594005};
test_output[3194] = '{0.193957847702};
############ END DEBUG ############*/
test_input[25560:25567] = '{32'h4218f8de, 32'h42823323, 32'h421ce07d, 32'h413416b9, 32'hc250e0ca, 32'h42841000, 32'hc20c7c1d, 32'h4226bb2a};
test_label[3195] = '{32'h413416b9};
test_output[3195] = '{32'h425c6e7a};
/*############ DEBUG ############
test_input[25560:25567] = '{38.2430336733, 65.0998770381, 39.2192281874, 11.2555472777, -52.21952245, 66.0312474712, -35.1212051655, 41.6827773281};
test_label[3195] = '{11.2555472777};
test_output[3195] = '{55.1078870978};
############ END DEBUG ############*/
test_input[25568:25575] = '{32'hc20b04f5, 32'h4281816e, 32'h424ac953, 32'hc1a60189, 32'hc2961e50, 32'h41aabbaf, 32'h41f69f02, 32'h42231ef3};
test_label[3196] = '{32'h42231ef3};
test_output[3196] = '{32'h41bfc7d4};
/*############ DEBUG ############
test_input[25568:25575] = '{-34.7548410095, 64.7527953982, 50.6966042933, -20.7507493487, -75.0592028918, 21.3416419603, 30.8276407237, 40.7802234475};
test_label[3196] = '{40.7802234475};
test_output[3196] = '{23.9725727368};
############ END DEBUG ############*/
test_input[25576:25583] = '{32'hc2935edf, 32'h42826498, 32'h42797e47, 32'h42027ad6, 32'hc21bb635, 32'hc215d75d, 32'hc291c112, 32'h424ca240};
test_label[3197] = '{32'hc2935edf};
test_output[3197] = '{32'h430af083};
/*############ DEBUG ############
test_input[25576:25583] = '{-73.685298029, 65.1964754689, 62.3733187055, 32.6199566065, -38.9279378263, -37.4603173807, -72.8770884673, 51.158449007};
test_label[3197] = '{-73.685298029};
test_output[3197] = '{138.939494027};
############ END DEBUG ############*/
test_input[25584:25591] = '{32'hc2b79e84, 32'h41aa8377, 32'hc2acd889, 32'h41ea0f3d, 32'h42c5de92, 32'hc2aa670a, 32'hc2a71848, 32'hc29e0682};
test_label[3198] = '{32'hc2acd889};
test_output[3198] = '{32'h43395b8e};
/*############ DEBUG ############
test_input[25584:25591] = '{-91.8095994936, 21.3141912663, -86.4229234381, 29.2574397939, 98.9347068724, -85.2012491727, -83.5474255292, -79.0127103963};
test_label[3198] = '{-86.4229234381};
test_output[3198] = '{185.35763031};
############ END DEBUG ############*/
test_input[25592:25599] = '{32'h41c315d5, 32'h420c4f46, 32'h3f3d069b, 32'hc2100c6b, 32'h42671735, 32'hc2020cbd, 32'hc2101f4e, 32'h427cb990};
test_label[3199] = '{32'h427cb990};
test_output[3199] = '{32'h3b926970};
/*############ DEBUG ############
test_input[25592:25599] = '{24.3856597184, 35.0774136387, 0.738382067536, -36.0121255173, 57.7726627497, -32.5124401269, -36.0305708026, 63.1812119251};
test_label[3199] = '{63.1812119251};
test_output[3199] = '{0.00446813548475};
############ END DEBUG ############*/
test_input[25600:25607] = '{32'hc27e6fa8, 32'hc1eda586, 32'h42b03280, 32'hc226a54b, 32'h425f4862, 32'hc201f362, 32'hc2650cc0, 32'hc1bf6093};
test_label[3200] = '{32'hc1eda586};
test_output[3200] = '{32'h42eb9be1};
/*############ DEBUG ############
test_input[25600:25607] = '{-63.6090394546, -29.7058215405, 88.0986290915, -41.661419762, 55.8206876461, -32.4876793462, -57.262450045, -23.9221554281};
test_label[3200] = '{-29.7058215405};
test_output[3200] = '{117.804450632};
############ END DEBUG ############*/
test_input[25608:25615] = '{32'hc17d0086, 32'hc27702de, 32'hc1ca3770, 32'h40572b01, 32'h42b30f24, 32'hc2c1f520, 32'hc2c503b5, 32'hc2c11f7a};
test_label[3201] = '{32'hc27702de};
test_output[3201] = '{32'h4317484a};
/*############ DEBUG ############
test_input[25608:25615] = '{-15.8126279355, -61.7528017489, -25.2770682354, 3.36199985259, 89.5295704587, -96.9787575075, -98.5072422746, -96.5614747933};
test_label[3201] = '{-61.7528017489};
test_output[3201] = '{151.282372208};
############ END DEBUG ############*/
test_input[25616:25623] = '{32'hc28cb9b0, 32'h429dcc02, 32'h41953682, 32'hc2a788ac, 32'hc2284f9c, 32'h41f1ede0, 32'hc2a26c70, 32'h41d9e2b4};
test_label[3202] = '{32'h41d9e2b4};
test_output[3202] = '{32'h424ea6ab};
/*############ DEBUG ############
test_input[25616:25623] = '{-70.3626729569, 78.8984564063, 18.6516149364, -83.7669387428, -42.0777416284, 30.2411492799, -81.2117911951, 27.2356950545};
test_label[3202] = '{27.2356950545};
test_output[3202] = '{51.6627613518};
############ END DEBUG ############*/
test_input[25624:25631] = '{32'h42068203, 32'hc1988a68, 32'hc22f0c0b, 32'h4238738e, 32'hc1921f80, 32'hc2abd480, 32'h428532d9, 32'hc1eb2336};
test_label[3203] = '{32'h428532d9};
test_output[3203] = '{32'h30ae297d};
/*############ DEBUG ############
test_input[25624:25631] = '{33.6269661547, -19.0675806151, -43.7617590473, 46.1128475371, -18.2653817315, -85.9150420872, 66.5993107653, -29.3921926924};
test_label[3203] = '{66.5993107653};
test_output[3203] = '{1.26719579355e-09};
############ END DEBUG ############*/
test_input[25632:25639] = '{32'hc1df7133, 32'h42b4db63, 32'hc1bbf83d, 32'h42342f4d, 32'hc20c07d2, 32'h40e75329, 32'hc0d4f567, 32'hc27be9d9};
test_label[3204] = '{32'hc1bbf83d};
test_output[3204] = '{32'h42e3d972};
/*############ DEBUG ############
test_input[25632:25639] = '{-27.930273783, 90.4284867869, -23.4962091852, 45.0461936759, -35.007637111, 7.22890141079, -6.65495641853, -62.9783670953};
test_label[3204] = '{-23.4962091852};
test_output[3204] = '{113.924695972};
############ END DEBUG ############*/
test_input[25640:25647] = '{32'h41b7c30c, 32'h42bc1c8d, 32'h41804038, 32'hc2a39883, 32'h419a20ca, 32'h41213ec7, 32'h4240a686, 32'hc2a9202d};
test_label[3205] = '{32'h4240a686};
test_output[3205] = '{32'h42379293};
/*############ DEBUG ############
test_input[25640:25647] = '{22.9702386096, 94.0557599743, 16.0313568607, -81.797876077, 19.266010056, 10.0778267019, 48.1626222706, -84.5628414522};
test_label[3205] = '{48.1626222706};
test_output[3205] = '{45.8931377036};
############ END DEBUG ############*/
test_input[25648:25655] = '{32'hc10769e6, 32'h424ce28e, 32'hc1814375, 32'hc24c3574, 32'hc17dc3c6, 32'hc20640f0, 32'hc2bf59b4, 32'hc221ca10};
test_label[3206] = '{32'hc20640f0};
test_output[3206] = '{32'h42a991bf};
/*############ DEBUG ############
test_input[25648:25655] = '{-8.46335363982, 51.2212455562, -16.1579381398, -51.0522020988, -15.8602967228, -33.5634171221, -95.6752001219, -40.447326887};
test_label[3206] = '{-33.5634171221};
test_output[3206] = '{84.7846626783};
############ END DEBUG ############*/
test_input[25656:25663] = '{32'hc2c46762, 32'h42b6adc4, 32'hc21eaf47, 32'h424ea6e3, 32'hc27060ab, 32'hc27dcea4, 32'h408afad6, 32'h4297f5b7};
test_label[3207] = '{32'h4297f5b7};
test_output[3207] = '{32'h4175c067};
/*############ DEBUG ############
test_input[25656:25663] = '{-98.2019207658, 91.33938302, -39.6711693481, 51.6629750543, -60.094403306, -63.4517985556, 4.34311976701, 75.979909786};
test_label[3207] = '{75.979909786};
test_output[3207] = '{15.3594734475};
############ END DEBUG ############*/
test_input[25664:25671] = '{32'h41d00a35, 32'hc14b4b6a, 32'hc197b45b, 32'h4261b524, 32'hc2638be0, 32'h4237f986, 32'h423748d5, 32'hc2ba4ccd};
test_label[3208] = '{32'hc197b45b};
test_output[3208] = '{32'h4296c7b0};
/*############ DEBUG ############
test_input[25664:25671] = '{26.0049841474, -12.7059119516, -18.963064004, 56.4268950385, -56.8865958788, 45.9936751323, 45.8211248732, -93.1499981576};
test_label[3208] = '{-18.963064004};
test_output[3208] = '{75.3900132518};
############ END DEBUG ############*/
test_input[25672:25679] = '{32'hc227ac0d, 32'h41d8c2d0, 32'h42a0f4f7, 32'hc1db2e45, 32'h42837a95, 32'h42be6220, 32'h40bc57b2, 32'hc2ade90a};
test_label[3209] = '{32'hc1db2e45};
test_output[3209] = '{32'h42f52db1};
/*############ DEBUG ############
test_input[25672:25679] = '{-41.9180170078, 27.0951240654, 80.4784449522, -27.3975928324, 65.7394197448, 95.1916511682, 5.88570491439, -86.9551538785};
test_label[3209] = '{-27.3975928324};
test_output[3209] = '{122.589244408};
############ END DEBUG ############*/
test_input[25680:25687] = '{32'h41c18474, 32'h424bb7ab, 32'hc28f4b50, 32'h42844680, 32'hc19a2543, 32'h42943125, 32'hc0b7be47, 32'h42b846dd};
test_label[3210] = '{32'h41c18474};
test_output[3210] = '{32'h4287e5c0};
/*############ DEBUG ############
test_input[25680:25687] = '{24.1896735918, 50.9293644819, -71.6470913061, 66.1376966812, -19.2681942356, 74.0959872879, -5.74197713217, 92.1384018475};
test_label[3210] = '{24.1896735918};
test_output[3210] = '{67.9487282703};
############ END DEBUG ############*/
test_input[25688:25695] = '{32'hc1a5b377, 32'h412fba74, 32'h4296a39e, 32'h420a8321, 32'hc23e2506, 32'h40a1d022, 32'hc0d8c76f, 32'h4296d073};
test_label[3211] = '{32'h420a8321};
test_output[3211] = '{32'h4225b7b4};
/*############ DEBUG ############
test_input[25688:25695] = '{-20.7126286622, 10.9830205, 75.319561607, 34.628054882, -47.5361549335, 5.05665689279, -6.77434483625, 75.4071299721};
test_label[3211] = '{34.628054882};
test_output[3211] = '{41.4293963093};
############ END DEBUG ############*/
test_input[25696:25703] = '{32'h42a6bfd2, 32'hc29d2197, 32'hc110bd03, 32'h41bdd143, 32'hc2324888, 32'h42929f3a, 32'hc2b6ce73, 32'hc272946c};
test_label[3212] = '{32'hc29d2197};
test_output[3212] = '{32'h4321f0b7};
/*############ DEBUG ############
test_input[25696:25703] = '{83.3746502357, -78.5656063422, -9.0461450938, 23.7271780803, -44.5708321692, 73.3109896107, -91.4032235943, -60.6449443694};
test_label[3212] = '{-78.5656063422};
test_output[3212] = '{161.940299177};
############ END DEBUG ############*/
test_input[25704:25711] = '{32'h418efce0, 32'hc2212e13, 32'hc23cd0ea, 32'hc1352b71, 32'h42a8ae7c, 32'hc0d08cb1, 32'h4217cf9f, 32'h42b9d62a};
test_label[3213] = '{32'hc23cd0ea};
test_output[3213] = '{32'h430c1f5c};
/*############ DEBUG ############
test_input[25704:25711] = '{17.8734744981, -40.2949927857, -47.2040161476, -11.3231060217, 84.34078785, -6.51717427123, 37.9527532012, 92.9182903775};
test_label[3213] = '{-47.2040161476};
test_output[3213] = '{140.122494802};
############ END DEBUG ############*/
test_input[25712:25719] = '{32'h4191c00d, 32'h419514c0, 32'h4207b1e6, 32'hc28f0273, 32'h421e10f1, 32'hc2bea890, 32'h42b9448c, 32'hc09f1966};
test_label[3214] = '{32'hc28f0273};
test_output[3214] = '{32'h4324237f};
/*############ DEBUG ############
test_input[25712:25719] = '{18.2187747595, 18.6351312959, 33.9237270953, -71.5047856724, 39.5165429048, -95.3292244071, 92.6338776475, -4.97185049647};
test_label[3214] = '{-71.5047856724};
test_output[3214] = '{164.13866332};
############ END DEBUG ############*/
test_input[25720:25727] = '{32'h41af5956, 32'h41aa405c, 32'hc2bb609c, 32'h42721852, 32'hc2c1c797, 32'h42b6fb20, 32'h403ea975, 32'h422ec412};
test_label[3215] = '{32'h42b6fb20};
test_output[3215] = '{32'h29208000};
/*############ DEBUG ############
test_input[25720:25727] = '{21.9186202441, 21.281426302, -93.6886885419, 60.523748784, -96.8898258453, 91.4904794299, 2.97909272787, 43.6914764515};
test_label[3215] = '{91.4904794299};
test_output[3215] = '{3.56381590905e-14};
############ END DEBUG ############*/
test_input[25728:25735] = '{32'hc10a3dcc, 32'hc22fa48e, 32'hc2b44790, 32'hc0688e54, 32'hc240c28c, 32'h42844425, 32'hbfb27a43, 32'hbfc31d7d};
test_label[3216] = '{32'hbfb27a43};
test_output[3216] = '{32'h42870e0f};
/*############ DEBUG ############
test_input[25728:25735] = '{-8.64008665828, -43.9106977293, -90.1397684689, -3.63368702755, -48.1899863385, 66.133098303, -1.3943560934, -1.52433744531};
test_label[3216] = '{-1.3943560934};
test_output[3216] = '{67.5274543964};
############ END DEBUG ############*/
test_input[25736:25743] = '{32'h41bbe948, 32'h423d463e, 32'hc203801d, 32'h4182f33c, 32'hc1e328d6, 32'h408de727, 32'h41232c6d, 32'hc23c1725};
test_label[3217] = '{32'h423d463e};
test_output[3217] = '{32'h2e4504e0};
/*############ DEBUG ############
test_input[25736:25743] = '{23.4889073356, 47.3185941115, -32.8751093806, 16.3687658614, -28.3949388349, 4.43446695876, 10.1983460025, -47.0226016059};
test_label[3217] = '{47.3185941115};
test_output[3217] = '{4.47969439331e-11};
############ END DEBUG ############*/
test_input[25744:25751] = '{32'hc20df31d, 32'hc18770cd, 32'h421390d7, 32'hc0a12f75, 32'hc28062cd, 32'h403cd7e8, 32'hc04fbbb9, 32'h429b43b7};
test_label[3218] = '{32'hc18770cd};
test_output[3218] = '{32'h42bd1fea};
/*############ DEBUG ############
test_input[25744:25751] = '{-35.4874170827, -16.9300776087, 36.8914469753, -5.03704314109, -64.1929701905, 2.95067791683, -3.24583262365, 77.6322530128};
test_label[3218] = '{-16.9300776087};
test_output[3218] = '{94.5623306215};
############ END DEBUG ############*/
test_input[25752:25759] = '{32'h429c7d91, 32'hc1a5ce14, 32'h429a6ffc, 32'hc24af049, 32'hc2a28da3, 32'h4168d537, 32'h42127e6d, 32'h4202eba9};
test_label[3219] = '{32'h429c7d91};
test_output[3219] = '{32'h3e9cc5b6};
/*############ DEBUG ############
test_input[25752:25759] = '{78.2452489006, -20.7256240738, 77.2187201399, -50.7346537425, -81.2766379553, 14.5520540068, 36.6234608497, 32.7301355299};
test_label[3219] = '{78.2452489006};
test_output[3219] = '{0.306195906768};
############ END DEBUG ############*/
test_input[25760:25767] = '{32'h42097a17, 32'h40844e96, 32'hc2811ad2, 32'h42be3ba1, 32'h427d3988, 32'h408385e9, 32'h4127fa9e, 32'hc2643ebe};
test_label[3220] = '{32'h42be3ba1};
test_output[3220] = '{32'h288b0000};
/*############ DEBUG ############
test_input[25760:25767] = '{34.3692279715, 4.1345927754, -64.5523800333, 95.116465177, 63.3061842254, 4.11009638335, 10.4986857586, -57.061271345};
test_label[3220] = '{95.116465177};
test_output[3220] = '{1.54321000423e-14};
############ END DEBUG ############*/
test_input[25768:25775] = '{32'h41ada9b2, 32'hc2c39b5e, 32'hc267905e, 32'hc23b9795, 32'hc2afb381, 32'h4230a91e, 32'hc1b8199b, 32'h426236e4};
test_label[3221] = '{32'h41ada9b2};
test_output[3221] = '{32'h420b620c};
/*############ DEBUG ############
test_input[25768:25775] = '{21.7078581493, -97.8034538, -57.8909819066, -46.8980282737, -87.8505973279, 44.1651543265, -23.0125023456, 56.5536043084};
test_label[3221] = '{21.7078581493};
test_output[3221] = '{34.8457503255};
############ END DEBUG ############*/
test_input[25776:25783] = '{32'hc2b040c7, 32'h42808e7e, 32'h42bebecf, 32'hc168d573, 32'h42afd3b2, 32'h42a91c3b, 32'hc15b00e2, 32'hbfbb8cee};
test_label[3222] = '{32'hc168d573};
test_output[3222] = '{32'h42dbd9cb};
/*############ DEBUG ############
test_input[25776:25783] = '{-88.1265170386, 64.2783053442, 95.37267329, -14.5521113817, 87.9134655151, 84.5551343671, -13.6877154755, -1.46523828414};
test_label[3222] = '{-14.5521113817};
test_output[3222] = '{109.925380651};
############ END DEBUG ############*/
test_input[25784:25791] = '{32'h41a86fb5, 32'h423fc4d5, 32'h428c3141, 32'hc2c770ef, 32'hc293ac3e, 32'hc2bf08f7, 32'hc2ab4e0e, 32'hc15a4a25};
test_label[3223] = '{32'hc2c770ef};
test_output[3223] = '{32'h4329d118};
/*############ DEBUG ############
test_input[25784:25791] = '{21.0545445781, 47.9422199594, 70.0961983393, -99.7205716667, -73.8364114762, -95.5175057807, -85.6524519616, -13.6431015805};
test_label[3223] = '{-99.7205716667};
test_output[3223] = '{169.816770006};
############ END DEBUG ############*/
test_input[25792:25799] = '{32'h428285f7, 32'hc1cee8db, 32'hc13a4701, 32'h422d2204, 32'h428b41f5, 32'hc2b58f38, 32'h425ceec8, 32'hc140bd3b};
test_label[3224] = '{32'hc140bd3b};
test_output[3224] = '{32'h42a36011};
/*############ DEBUG ############
test_input[25792:25799] = '{65.2616463024, -25.8636986801, -11.6423346727, 43.2832198999, 69.6288239358, -90.7797247354, 55.2331832272, -12.0461985218};
test_label[3224] = '{-12.0461985218};
test_output[3224] = '{81.6876302022};
############ END DEBUG ############*/
test_input[25800:25807] = '{32'hc24736f6, 32'h418b1f5e, 32'h42c6b61a, 32'hc19656e9, 32'hc2abd5e8, 32'hc11626ac, 32'h4249c9e6, 32'hc22e3a3b};
test_label[3225] = '{32'hc22e3a3b};
test_output[3225] = '{32'h430ee99c};
/*############ DEBUG ############
test_input[25800:25807] = '{-49.8036719863, 17.3903162406, 99.3556642347, -18.7924368292, -85.9177851703, -9.38444176355, 50.4471683087, -43.5568647833};
test_label[3225] = '{-43.5568647833};
test_output[3225] = '{142.912529018};
############ END DEBUG ############*/
test_input[25808:25815] = '{32'h42253992, 32'h41e6090b, 32'hc1ec55f1, 32'hc288eb9e, 32'h4259967b, 32'h428a8581, 32'h426ca4e7, 32'hc2ba23a0};
test_label[3226] = '{32'hc2ba23a0};
test_output[3226] = '{32'h43225493};
/*############ DEBUG ############
test_input[25808:25815] = '{41.306220747, 28.7544158808, -29.5419638422, -68.4601879242, 54.3969524494, 69.2607465785, 59.1610387452, -93.0695784742};
test_label[3226] = '{-93.0695784742};
test_output[3226] = '{162.330366494};
############ END DEBUG ############*/
test_input[25816:25823] = '{32'hc291d0f3, 32'hc1819492, 32'hc291d7da, 32'hc16c58bc, 32'hc2007f14, 32'h428f4015, 32'h4292f5ee, 32'hc2ac6a65};
test_label[3227] = '{32'hc16c58bc};
test_output[3227] = '{32'h42b0cb6f};
/*############ DEBUG ############
test_input[25816:25823] = '{-72.9081072171, -16.1975438269, -72.9215877625, -14.7716634605, -32.1240982031, 71.6251593737, 73.4803310221, -86.2078030462};
test_label[3227] = '{-14.7716634605};
test_output[3227] = '{88.397328775};
############ END DEBUG ############*/
test_input[25824:25831] = '{32'h4210b230, 32'hc209df0b, 32'hc28981fc, 32'h4228be1f, 32'h41945ba0, 32'hc256c16d, 32'h3f92fa18, 32'hc1bde059};
test_label[3228] = '{32'h4228be1f};
test_output[3228] = '{32'h3b205e72};
/*############ DEBUG ############
test_input[25824:25831] = '{36.1740116578, -34.4678143412, -68.7538756948, 42.1856658266, 18.5447380575, -53.6888915012, 1.14825730898, -23.7345451678};
test_label[3228] = '{42.1856658266};
test_output[3228] = '{0.00244703567865};
############ END DEBUG ############*/
test_input[25832:25839] = '{32'hc24229b9, 32'h426637ac, 32'hc211884e, 32'hc23ade0b, 32'hc280dbc6, 32'hc20450ef, 32'hc16b0d1e, 32'hc1d5d375};
test_label[3229] = '{32'hc20450ef};
test_output[3229] = '{32'h42b5444d};
/*############ DEBUG ############
test_input[25832:25839] = '{-48.5407435802, 57.5543652274, -36.3831083612, -46.7168399028, -64.4292482863, -33.0790370501, -14.6907026124, -26.7282498557};
test_label[3229] = '{-33.0790370501};
test_output[3229] = '{90.6334022775};
############ END DEBUG ############*/
test_input[25840:25847] = '{32'h42a95bda, 32'h41a21c03, 32'h4067635b, 32'h4291db4b, 32'hc1d581bf, 32'hc0cca78c, 32'h41494731, 32'h429822b7};
test_label[3230] = '{32'hc1d581bf};
test_output[3230] = '{32'h42debc63};
/*############ DEBUG ############
test_input[25840:25847] = '{84.6793971759, 20.263678472, 3.61543916325, 72.9283089347, -26.6883525597, -6.39545265738, 12.579880732, 76.0678054141};
test_label[3230] = '{-26.6883525597};
test_output[3230] = '{111.367939582};
############ END DEBUG ############*/
test_input[25848:25855] = '{32'hc285ad92, 32'hc1b5aa64, 32'hc2be9bb7, 32'hc2936eb2, 32'h4288e65a, 32'h41f4a816, 32'h42be055d, 32'hc1adab2b};
test_label[3231] = '{32'h4288e65a};
test_output[3231] = '{32'h41d47c0c};
/*############ DEBUG ############
test_input[25848:25855] = '{-66.8390008175, -22.7081977598, -95.304128106, -73.7162011016, 68.4499071011, 30.5820727869, 95.0104765036, -21.7085776279};
test_label[3231] = '{68.4499071011};
test_output[3231] = '{26.5605694026};
############ END DEBUG ############*/
test_input[25856:25863] = '{32'h42362769, 32'hc2c5e870, 32'hc2258a5e, 32'hc21a4474, 32'h42808cec, 32'h425998e0, 32'h4105d57d, 32'hc24d2794};
test_label[3232] = '{32'hc21a4474};
test_output[3232] = '{32'h42cdaf2c};
/*############ DEBUG ############
test_input[25856:25863] = '{45.538487997, -98.9539823939, -41.3851254247, -38.5668483108, 64.2752365082, 54.399290708, 8.36462142819, -51.2886519362};
test_label[3232] = '{-38.5668483108};
test_output[3232] = '{102.842136221};
############ END DEBUG ############*/
test_input[25864:25871] = '{32'hc2aa6032, 32'h41be5f20, 32'hc1108a63, 32'h42a1ae9c, 32'h3f311564, 32'hc258d056, 32'h429b9921, 32'h41a2040c};
test_label[3233] = '{32'h41be5f20};
test_output[3233] = '{32'h42645d6b};
/*############ DEBUG ############
test_input[25864:25871] = '{-85.187880664, 23.7964468982, -9.03378614799, 80.8410372054, 0.691732636848, -54.2034522105, 77.7990802416, 20.2519758219};
test_label[3233] = '{23.7964468982};
test_output[3233] = '{57.0912270782};
############ END DEBUG ############*/
test_input[25872:25879] = '{32'hc2098ad5, 32'h4191a52e, 32'hc2b12b19, 32'hc25b0de3, 32'h42bd71b0, 32'hc26a296c, 32'hc2c25e3f, 32'hc2223a6e};
test_label[3234] = '{32'h42bd71b0};
test_output[3234] = '{32'h80000000};
/*############ DEBUG ############
test_input[25872:25879] = '{-34.3855792417, 18.2056535227, -88.5841772495, -54.7635627886, 94.7220491667, -58.5404510418, -97.1840768684, -40.5570601633};
test_label[3234] = '{94.7220491667};
test_output[3234] = '{-0.0};
############ END DEBUG ############*/
test_input[25880:25887] = '{32'h3ea43eb6, 32'h42ac1371, 32'hc1b7a331, 32'hc1f817d2, 32'hc26337bb, 32'h41d028b1, 32'hc12294ea, 32'hc2b61bb2};
test_label[3235] = '{32'h41d028b1};
test_output[3235] = '{32'h42701289};
/*############ DEBUG ############
test_input[25880:25887] = '{0.320790955797, 86.0379705193, -22.9546839163, -31.0116302272, -56.8044252374, 26.01986899, -10.161355782, -91.0540920049};
test_label[3235] = '{26.01986899};
test_output[3235] = '{60.0181015293};
############ END DEBUG ############*/
test_input[25888:25895] = '{32'hc2824a7b, 32'hc26569f5, 32'hc2392921, 32'h4250f044, 32'hc0635a8e, 32'hc1cadf33, 32'h42ba4831, 32'h40c43999};
test_label[3236] = '{32'hc1cadf33};
test_output[3236] = '{32'h42ecfffe};
/*############ DEBUG ############
test_input[25888:25895] = '{-65.1454730901, -57.3534755025, -46.2901651291, 52.2346358195, -3.55240194127, -25.3589841336, 93.1409971945, 6.13203076883};
test_label[3236] = '{-25.3589841336};
test_output[3236] = '{118.499981328};
############ END DEBUG ############*/
test_input[25896:25903] = '{32'h3e494e74, 32'h4234f834, 32'hc1773a01, 32'h422f4e61, 32'hc2c0675d, 32'hc1512cb0, 32'h41bc55d0, 32'h4218c098};
test_label[3237] = '{32'hc2c0675d};
test_output[3237] = '{32'h430da98a};
/*############ DEBUG ############
test_input[25896:25903] = '{0.196588334298, 45.2423868649, -15.4516611336, 43.8265418014, -96.201884151, -13.07340958, 23.5419012419, 38.1880780543};
test_label[3237] = '{-96.201884151};
test_output[3237] = '{141.662268624};
############ END DEBUG ############*/
test_input[25904:25911] = '{32'h4285e865, 32'h4291cfa1, 32'h42278c20, 32'h41aa9191, 32'h429a1916, 32'hc2731b5b, 32'hc21f55f3, 32'h42368b65};
test_label[3238] = '{32'h42278c20};
test_output[3238] = '{32'h420cb636};
/*############ DEBUG ############
test_input[25904:25911] = '{66.9538970118, 72.9055262342, 41.8868398224, 21.3210767638, 77.0489983334, -60.7767136815, -39.8339350394, 45.6361289687};
test_label[3238] = '{41.8868398224};
test_output[3238] = '{35.177942233};
############ END DEBUG ############*/
test_input[25912:25919] = '{32'h42b62c42, 32'hc19f9654, 32'hc25d4827, 32'h41a093af, 32'h421f880e, 32'h4237b295, 32'h421509f6, 32'h42c2e712};
test_label[3239] = '{32'h421f880e};
test_output[3239] = '{32'h426647d8};
/*############ DEBUG ############
test_input[25912:25919] = '{91.0864416021, -19.9484020933, -55.3204610865, 20.0721107549, 39.8828665808, 45.9243953098, 37.2597283558, 97.4513074501};
test_label[3239] = '{39.8828665808};
test_output[3239] = '{57.5701603624};
############ END DEBUG ############*/
test_input[25920:25927] = '{32'hc29e645a, 32'hc23aa476, 32'h429c44dc, 32'hc1db7682, 32'h4211fb86, 32'h420f7034, 32'hc16097d7, 32'h41a074da};
test_label[3240] = '{32'hc16097d7};
test_output[3240] = '{32'h42b857d7};
/*############ DEBUG ############
test_input[25920:25927] = '{-79.1959989841, -46.6606056217, 78.1344920513, -27.432864575, 36.4956287724, 35.8595735021, -14.0370703713, 20.0570560929};
test_label[3240] = '{-14.0370703713};
test_output[3240] = '{92.1715624226};
############ END DEBUG ############*/
test_input[25928:25935] = '{32'h40f7bdc9, 32'hc01679dd, 32'h421dffc9, 32'h42ad0a52, 32'hc2a9737b, 32'hc2b5f2e7, 32'hc1e943d8, 32'hc2bed2d7};
test_label[3241] = '{32'hc2a9737b};
test_output[3241] = '{32'h432b3ee7};
/*############ DEBUG ############
test_input[25928:25935] = '{7.74191705753, -2.35118787861, 39.4997908189, 86.5201580946, -84.7255486635, -90.9744212411, -29.158126309, -95.4117959837};
test_label[3241] = '{-84.7255486635};
test_output[3241] = '{171.245706758};
############ END DEBUG ############*/
test_input[25936:25943] = '{32'h4216b082, 32'h42acbd31, 32'hc2a0d2a3, 32'hc2a9c550, 32'h42c3bcbf, 32'h42ba80b0, 32'h42390a2b, 32'hc2c0172a};
test_label[3242] = '{32'hc2c0172a};
test_output[3242] = '{32'h4341ec7a};
/*############ DEBUG ############
test_input[25936:25943] = '{37.6723697249, 86.3695108983, -80.4114029545, -84.8853782468, 97.8686482879, 93.2513454466, 46.2599293544, -96.0452460246};
test_label[3242] = '{-96.0452460246};
test_output[3242] = '{193.923735276};
############ END DEBUG ############*/
test_input[25944:25951] = '{32'hc2468602, 32'hc20a29b3, 32'hc1fb473d, 32'h41f40eae, 32'h4291a518, 32'hc238041a, 32'hc280a37f, 32'hc26569b9};
test_label[3243] = '{32'hc20a29b3};
test_output[3243] = '{32'h42d6b9f2};
/*############ DEBUG ############
test_input[25944:25951] = '{-49.6308685233, -34.5407214829, -31.4097849952, 30.5071685085, 72.8224495354, -46.0040042768, -64.319331513, -57.3532437378};
test_label[3243] = '{-34.5407214829};
test_output[3243] = '{107.363171018};
############ END DEBUG ############*/
test_input[25952:25959] = '{32'h422acb87, 32'hc1e96ef1, 32'h42683cec, 32'h4282c6d3, 32'h41e555b8, 32'hc23c0a5b, 32'hc2b13878, 32'h42c4317c};
test_label[3244] = '{32'hc23c0a5b};
test_output[3244] = '{32'h43111b55};
/*############ DEBUG ############
test_input[25952:25959] = '{42.698759004, -29.1791707893, 58.0594933494, 65.3883258316, 28.6668546267, -47.0101112569, -88.6102906779, 98.0966500186};
test_label[3244] = '{-47.0101112569};
test_output[3244] = '{145.106761276};
############ END DEBUG ############*/
test_input[25960:25967] = '{32'h42b52217, 32'h40b7cc3c, 32'h42835abc, 32'h41ed1d98, 32'hc2a61688, 32'h42aabf43, 32'h42523a0a, 32'h42ab82a0};
test_label[3245] = '{32'h41ed1d98};
test_output[3245] = '{32'h4273c34e};
/*############ DEBUG ############
test_input[25960:25967] = '{90.5665799301, 5.74368090153, 65.6772143576, 29.6394500346, -83.0440066417, 85.3735618124, 52.5566804266, 85.7551264443};
test_label[3245] = '{29.6394500346};
test_output[3245] = '{60.940728258};
############ END DEBUG ############*/
test_input[25968:25975] = '{32'hc1a0e254, 32'h42b3b09d, 32'h42a89b46, 32'h42540dd3, 32'hc2288981, 32'hc1ce3959, 32'h40e91a34, 32'h42702d76};
test_label[3246] = '{32'hc1a0e254};
test_output[3246] = '{32'h42dbeb33};
/*############ DEBUG ############
test_input[25968:25975] = '{-20.1105108331, 89.8449499186, 84.3032646734, 53.0135010013, -42.1342797745, -25.77800102, 7.28444871007, 60.0443939812};
test_label[3246] = '{-20.1105108331};
test_output[3246] = '{109.959373004};
############ END DEBUG ############*/
test_input[25976:25983] = '{32'h42c3df16, 32'hc22e5088, 32'h42c3d902, 32'h41379d8e, 32'hc178dc21, 32'h42980ea5, 32'h41e16ec6, 32'hc270b691};
test_label[3247] = '{32'hc270b691};
test_output[3247] = '{32'h431ecd1e};
/*############ DEBUG ############
test_input[25976:25983] = '{97.9357170397, -43.5786448976, 97.9238445525, 11.4759658265, -15.5537428337, 76.0285995575, 28.1790890891, -60.1782886777};
test_label[3247] = '{-60.1782886777};
test_output[3247] = '{158.801234274};
############ END DEBUG ############*/
test_input[25984:25991] = '{32'hc2981abe, 32'h4199f4c3, 32'h40d90293, 32'h40a4af63, 32'hc1f7ddcb, 32'h424ff862, 32'hc29f213a, 32'hc18b16ad};
test_label[3248] = '{32'h424ff862};
test_output[3248] = '{32'h27d80000};
/*############ DEBUG ############
test_input[25984:25991] = '{-76.0522279787, 19.2445126642, 6.7815641962, 5.14640944958, -30.9832981292, 51.9925602922, -79.5648929848, -17.3860726052};
test_label[3248] = '{51.9925602922};
test_output[3248] = '{5.99520433298e-15};
############ END DEBUG ############*/
test_input[25992:25999] = '{32'h40490558, 32'hc29d1332, 32'h42a2f645, 32'hc17d3a95, 32'h417cf8c5, 32'h4219366c, 32'hbf9e8c2b, 32'h42a8e403};
test_label[3249] = '{32'hbf9e8c2b};
test_output[3249] = '{32'h42ab77f5};
/*############ DEBUG ############
test_input[25992:25999] = '{3.14095111423, -78.5374892231, 81.4809969406, -15.8268018997, 15.8107345968, 38.3031469571, -1.2386526394, 84.4453321985};
test_label[3249] = '{-1.2386526394};
test_output[3249] = '{85.7342926642};
############ END DEBUG ############*/
test_input[26000:26007] = '{32'h42b9f719, 32'hc23e466a, 32'hc2a28f51, 32'h42b2d3c5, 32'hc27e2837, 32'h4295f42a, 32'hc1af44e9, 32'h4293c123};
test_label[3250] = '{32'hc23e466a};
test_output[3250] = '{32'h430c9444};
/*############ DEBUG ############
test_input[26000:26007] = '{92.9826112198, -47.5687636142, -81.2799142925, 89.4136142946, -63.539270945, 74.9768863995, -21.9086466908, 73.8772171699};
test_label[3250] = '{-47.5687636142};
test_output[3250] = '{140.5791691};
############ END DEBUG ############*/
test_input[26008:26015] = '{32'h42a55921, 32'h42a638b0, 32'hc2bf3ec4, 32'hc1cb4b3f, 32'h4297948a, 32'hc12e9188, 32'h429107cd, 32'h4285e533};
test_label[3251] = '{32'h429107cd};
test_output[3251] = '{32'h4131828f};
/*############ DEBUG ############
test_input[26008:26015] = '{82.6740784599, 83.1107179864, -95.6225872733, -25.4117409485, 75.7901134759, -10.9105303299, 72.5152328805, 66.9476566635};
test_label[3251] = '{72.5152328805};
test_output[3251] = '{11.0943745047};
############ END DEBUG ############*/
test_input[26016:26023] = '{32'h4280f031, 32'hc2598720, 32'h415a0968, 32'h42762746, 32'h4291471a, 32'h41ddea60, 32'hc1b0ab33, 32'h4159e5ab};
test_label[3252] = '{32'h415a0968};
test_output[3252] = '{32'h426c0c28};
/*############ DEBUG ############
test_input[26016:26023] = '{64.469125437, -54.3819575156, 13.6272966725, 61.5383545346, 72.6388714226, 27.7394410585, -22.0835941623, 13.6185708057};
test_label[3252] = '{13.6272966725};
test_output[3252] = '{59.0118729001};
############ END DEBUG ############*/
test_input[26024:26031] = '{32'h42904d87, 32'h42a7868f, 32'h42afef7d, 32'h42b20d6c, 32'hc19a0c28, 32'h4298b63c, 32'hc2136b19, 32'h42149e56};
test_label[3253] = '{32'h42afef7d};
test_output[3253] = '{32'h3fae1a26};
/*############ DEBUG ############
test_input[26024:26031] = '{72.1514193082, 83.7628115024, 87.9677491299, 89.0262115759, -19.2559352722, 76.3559272015, -36.8545889097, 37.1546266003};
test_label[3253] = '{87.9677491299};
test_output[3253] = '{1.36017298892};
############ END DEBUG ############*/
test_input[26032:26039] = '{32'h41ea3bdb, 32'hc242f47a, 32'h419f2688, 32'h4201c5ba, 32'hc1942176, 32'hc29d9e73, 32'hc182c853, 32'hc29aa07f};
test_label[3254] = '{32'hc29d9e73};
test_output[3254] = '{32'h42de9682};
/*############ DEBUG ############
test_input[26032:26039] = '{29.2792263659, -48.7387449729, 19.8938135383, 32.4430919701, -18.5163388927, -78.8094721042, -16.3478145718, -77.3134656374};
test_label[3254] = '{-78.8094721042};
test_output[3254] = '{111.293960883};
############ END DEBUG ############*/
test_input[26040:26047] = '{32'h42b139f2, 32'hc2a11c04, 32'hc2817497, 32'h41af3e25, 32'hc125a4d0, 32'hc2402683, 32'hc2b4e2a8, 32'h421e1a1e};
test_label[3255] = '{32'h42b139f2};
test_output[3255] = '{32'h80000000};
/*############ DEBUG ############
test_input[26040:26047] = '{88.6131748655, -80.554716283, -64.7277147941, 21.9053445335, -10.3527376818, -48.0376091875, -90.4426874236, 39.5255057134};
test_label[3255] = '{88.6131748655};
test_output[3255] = '{-0.0};
############ END DEBUG ############*/
test_input[26048:26055] = '{32'hc219d1b5, 32'h42631895, 32'h428b41a1, 32'hc23f73bc, 32'hc10247f7, 32'hc164b746, 32'h42526984, 32'h426d940f};
test_label[3256] = '{32'h428b41a1};
test_output[3256] = '{32'h3821e365};
/*############ DEBUG ############
test_input[26048:26055] = '{-38.4547903717, 56.7740071404, 69.6281839167, -47.863020488, -8.1425695032, -14.2947443529, 52.6030443614, 59.3945899369};
test_label[3256] = '{69.6281839167};
test_output[3256] = '{3.85971701589e-05};
############ END DEBUG ############*/
test_input[26056:26063] = '{32'hc188678c, 32'hc29f70e4, 32'hc0d4e0ee, 32'h40755da8, 32'hc2932da9, 32'hc1bb2068, 32'hc2c5b347, 32'h4185ac07};
test_label[3257] = '{32'hc1bb2068};
test_output[3257] = '{32'h42206638};
/*############ DEBUG ############
test_input[26056:26063] = '{-17.0505607348, -79.7204905721, -6.65245746375, 3.83384121718, -73.5891802658, -23.3908242964, -98.8501526023, 16.7089976021};
test_label[3257] = '{-23.3908242964};
test_output[3257] = '{40.0998244594};
############ END DEBUG ############*/
test_input[26064:26071] = '{32'hc200c2f7, 32'h427813b6, 32'h4286c20e, 32'h42a42776, 32'h428ef6fe, 32'hc29a07d6, 32'h4184e895, 32'hc293ad38};
test_label[3258] = '{32'h4286c20e};
test_output[3258] = '{32'h416b2b62};
/*############ DEBUG ############
test_input[26064:26071] = '{-32.1903941885, 62.0192473287, 67.3790093747, 82.0770754936, 71.4824070726, -77.0153064491, 16.6135657299, -73.8383141871};
test_label[3258] = '{67.3790093747};
test_output[3258] = '{14.6980915835};
############ END DEBUG ############*/
test_input[26072:26079] = '{32'h4256577a, 32'hc2a24d85, 32'h4210e148, 32'h424a308a, 32'h41416b36, 32'hc2a6da6b, 32'hc14b6aa5, 32'hc2c62296};
test_label[3259] = '{32'h4256577a};
test_output[3259] = '{32'h3d3fc283};
/*############ DEBUG ############
test_input[26072:26079] = '{53.5854262565, -81.1514035133, 36.2200027221, 50.5474026327, 12.0886745701, -83.4265979854, -12.713535824, -99.067554215};
test_label[3259] = '{53.5854262565};
test_output[3259] = '{0.0468163617346};
############ END DEBUG ############*/
test_input[26080:26087] = '{32'h42bb411d, 32'hc2bf0e1a, 32'h41fb9d39, 32'hc1f8cb07, 32'h41cf4438, 32'hc29f67a0, 32'h42b95533, 32'h426c6521};
test_label[3260] = '{32'h42bb411d};
test_output[3260] = '{32'h3ea5ded9};
/*############ DEBUG ############
test_input[26080:26087] = '{93.6271722675, -95.5275386054, 31.4517688516, -31.0991353626, 25.9083101141, -79.7023936961, 92.6664071892, 59.0987595568};
test_label[3260] = '{93.6271722675};
test_output[3260] = '{0.323965824263};
############ END DEBUG ############*/
test_input[26088:26095] = '{32'hc12ec926, 32'h4235c559, 32'h42890edc, 32'hc2b6dd16, 32'hc2998d33, 32'h4296ba2f, 32'h420535b6, 32'h42170c6d};
test_label[3261] = '{32'h42890edc};
test_output[3261] = '{32'h40dabdf9};
/*############ DEBUG ############
test_input[26088:26095] = '{-10.9241083251, 45.4427213031, 68.5290212882, -91.4318086833, -76.7757808646, 75.3636360775, 33.302452762, 37.7621347219};
test_label[3261] = '{68.5290212882};
test_output[3261] = '{6.83569009265};
############ END DEBUG ############*/
test_input[26096:26103] = '{32'h4275a077, 32'hc17cbb70, 32'hc2476314, 32'hc0f551e4, 32'hc22f5721, 32'hc2a0c1cc, 32'hc2b999f8, 32'h42329dc7};
test_label[3262] = '{32'h42329dc7};
test_output[3262] = '{32'h41860560};
/*############ DEBUG ############
test_input[26096:26103] = '{61.4067053886, -15.7957610141, -49.8467573788, -7.66624664774, -43.8350886145, -80.3785094851, -92.8007216026, 44.6540804906};
test_label[3262] = '{44.6540804906};
test_output[3262] = '{16.7526249511};
############ END DEBUG ############*/
test_input[26104:26111] = '{32'h42789098, 32'h42397dd1, 32'hc23b70b1, 32'h427d9c65, 32'h40cde5fd, 32'h419a92f6, 32'hc2660196, 32'hc2ad854e};
test_label[3263] = '{32'h40cde5fd};
test_output[3263] = '{32'h4264df01};
/*############ DEBUG ############
test_input[26104:26111] = '{62.1412036104, 46.3728661174, -46.8600507502, 63.4027289211, 6.43432496159, 19.3217588045, -57.5015496812, -86.760363257};
test_label[3263] = '{6.43432496159};
test_output[3263] = '{57.2177778564};
############ END DEBUG ############*/
test_input[26112:26119] = '{32'hc2507981, 32'hc2b63474, 32'hc251fceb, 32'h429994d3, 32'hc1af0825, 32'h3ffee46e, 32'h42c5f000, 32'h424f8430};
test_label[3264] = '{32'hc251fceb};
test_output[3264] = '{32'h4317773b};
/*############ DEBUG ############
test_input[26112:26119] = '{-52.1186549915, -91.1024472779, -52.4969911909, 76.7906696362, -21.8789768567, 1.99134617838, 98.9687529192, 51.8790878694};
test_label[3264] = '{-52.4969911909};
test_output[3264] = '{151.46574411};
############ END DEBUG ############*/
test_input[26120:26127] = '{32'h423670cc, 32'hc290c1ce, 32'hc2a51d53, 32'h42276dcd, 32'hc277a5e4, 32'h42b17af5, 32'hc20872a7, 32'h4167c0aa};
test_label[3265] = '{32'h423670cc};
test_output[3265] = '{32'h422c851d};
/*############ DEBUG ############
test_input[26120:26127] = '{45.6101537675, -72.3785246489, -82.5572712791, 41.8572265513, -61.9120030683, 88.7401467513, -34.1119637752, 14.4845369421};
test_label[3265] = '{45.6101537675};
test_output[3265] = '{43.1299929838};
############ END DEBUG ############*/
test_input[26128:26135] = '{32'hc2c5dabe, 32'h4197ec4d, 32'h422bf609, 32'hc1d335b8, 32'h42b88464, 32'h42af6389, 32'h42ab25a1, 32'h42469375};
test_label[3266] = '{32'h42469375};
test_output[3266] = '{32'h422a8134};
/*############ DEBUG ############
test_input[26128:26135] = '{-98.9272323465, 18.9903817287, 42.9902695336, -26.4012298971, 92.2585754008, 87.6944067961, 85.573495626, 49.6440005789};
test_label[3266] = '{49.6440005789};
test_output[3266] = '{42.6261752288};
############ END DEBUG ############*/
test_input[26136:26143] = '{32'h4231c42f, 32'h428d4923, 32'hc243ff1a, 32'hc2b02603, 32'h42c4f546, 32'h428eaef6, 32'hc23cca4f, 32'h427db591};
test_label[3267] = '{32'h4231c42f};
test_output[3267] = '{32'h4258265d};
/*############ DEBUG ############
test_input[26136:26143] = '{44.4415866097, 70.6428481373, -48.9991228211, -88.0742381834, 98.4790489916, 71.3417181457, -47.1975685533, 63.4273091697};
test_label[3267] = '{44.4415866097};
test_output[3267] = '{54.0374623819};
############ END DEBUG ############*/
test_input[26144:26151] = '{32'hc23166ea, 32'hc0a36604, 32'hc28671d1, 32'hc2460454, 32'h41cde88e, 32'hc1f944ef, 32'h4182d0ed, 32'h42af6748};
test_label[3268] = '{32'hc2460454};
test_output[3268] = '{32'h430934b9};
/*############ DEBUG ############
test_input[26144:26151] = '{-44.3505015562, -5.10620302755, -67.2223007723, -49.5042250036, 25.7385513613, -31.1586590599, 16.3520147684, 87.7017181806};
test_label[3268] = '{-49.5042250036};
test_output[3268] = '{137.205943184};
############ END DEBUG ############*/
test_input[26152:26159] = '{32'h4170d82b, 32'h42c0e92b, 32'hc1095f44, 32'hc2951568, 32'hc05c7b5f, 32'h41eac97b, 32'h3e9548ad, 32'hc18cdf39};
test_label[3269] = '{32'hc1095f44};
test_output[3269] = '{32'h42d21513};
/*############ DEBUG ############
test_input[26152:26159] = '{15.0527752946, 96.4554031936, -8.58575778076, -74.5418058669, -3.44503004848, 29.348379262, 0.291570088087, -17.6089948075};
test_label[3269] = '{-8.58575778076};
test_output[3269] = '{105.041160974};
############ END DEBUG ############*/
test_input[26160:26167] = '{32'hc2bad36b, 32'hc25fa4f6, 32'hc24c4231, 32'hc240561e, 32'h4211ccb3, 32'h42424436, 32'h42af44ad, 32'hc2932c1e};
test_label[3270] = '{32'h42424436};
test_output[3270] = '{32'h421c4523};
/*############ DEBUG ############
test_input[26160:26167] = '{-93.4129255093, -55.9110961306, -51.0646381923, -48.0840969665, 36.4499013158, 48.5666121218, 87.63412938, -73.5861669515};
test_label[3270] = '{48.5666121218};
test_output[3270] = '{39.0675172582};
############ END DEBUG ############*/
test_input[26168:26175] = '{32'hc1e4e144, 32'hc2136066, 32'hc2ba6468, 32'hc293b737, 32'h40a19745, 32'h415d4a04, 32'h42b1a424, 32'hc2bc6164};
test_label[3271] = '{32'h42b1a424};
test_output[3271] = '{32'h80000000};
/*############ DEBUG ############
test_input[26168:26175] = '{-28.609992792, -36.8441382393, -93.1961035264, -73.8578415233, 5.04971554762, 13.8305699023, 88.820583937, -94.1902122972};
test_label[3271] = '{88.820583937};
test_output[3271] = '{-0.0};
############ END DEBUG ############*/
test_input[26176:26183] = '{32'h423a7a64, 32'h42b90161, 32'h42b666f0, 32'hc1c36047, 32'hc2a2f925, 32'h42b8fd22, 32'hc1b8c37f, 32'hc26cc076};
test_label[3272] = '{32'hc1c36047};
test_output[3272] = '{32'h42eb7bc8};
/*############ DEBUG ############
test_input[26176:26183] = '{46.6195231904, 92.5026906559, 91.2010523519, -24.4220102687, -81.4866086439, 92.49439637, -23.0954572316, -59.187951443};
test_label[3272] = '{-24.4220102687};
test_output[3272] = '{117.741757088};
############ END DEBUG ############*/
test_input[26184:26191] = '{32'hc18f2a3c, 32'hc25b7eff, 32'h42c65964, 32'hc2c435d8, 32'hc1429b75, 32'h42700121, 32'hc22dbf04, 32'h41f4e808};
test_label[3273] = '{32'hc1429b75};
test_output[3273] = '{32'h42deacd2};
/*############ DEBUG ############
test_input[26184:26191] = '{-17.8956218096, -54.8740189098, 99.1745877943, -98.1051638625, -12.162953032, 60.0011012342, -43.436538353, 30.6132960185};
test_label[3273] = '{-12.162953032};
test_output[3273] = '{111.337540826};
############ END DEBUG ############*/
test_input[26192:26199] = '{32'hc2b01ed0, 32'h42bcb129, 32'h42ab8516, 32'h421e286c, 32'hc1d57453, 32'hc1b04255, 32'hc21c4792, 32'hc1b28888};
test_label[3274] = '{32'h42ab8516};
test_output[3274] = '{32'h4109615f};
/*############ DEBUG ############
test_input[26192:26199] = '{-88.060182023, 94.3460191316, 85.7599333669, 39.5394730977, -26.681798952, -22.0323881525, -39.0698912245, -22.3166664887};
test_label[3274] = '{85.7599333669};
test_output[3274] = '{8.58627243273};
############ END DEBUG ############*/
test_input[26200:26207] = '{32'hc1876eec, 32'h4252ba46, 32'hc2ae44f2, 32'hc298fa9e, 32'h424c5019, 32'hc257d3fd, 32'hbfcd1f0e, 32'hc29a5079};
test_label[3275] = '{32'hc2ae44f2};
test_output[3275] = '{32'h430bfff6};
/*############ DEBUG ############
test_input[26200:26207] = '{-16.9291616481, 52.6819074676, -87.1346611935, -76.4894843841, 51.0782216515, -53.9570203638, -1.60251018896, -77.1571695589};
test_label[3275] = '{-87.1346611935};
test_output[3275] = '{139.999851201};
############ END DEBUG ############*/
test_input[26208:26215] = '{32'hc1412d2a, 32'hc086cc44, 32'h41b9d2b1, 32'h41688869, 32'hc2c224a2, 32'h422fa6ef, 32'hc280dd19, 32'hc2389113};
test_label[3276] = '{32'h41688869};
test_output[3276] = '{32'h41eb09aa};
/*############ DEBUG ############
test_input[26208:26215] = '{-12.073526746, -4.21243462599, 23.227876029, 14.5333035672, -97.0715482183, 43.9130229814, -64.4318285675, -46.1416757766};
test_label[3276] = '{14.5333035672};
test_output[3276] = '{29.3797194152};
############ END DEBUG ############*/
test_input[26216:26223] = '{32'hc2bb7a58, 32'hc20124e9, 32'hc272daf1, 32'h4267b9b2, 32'hc2aee6cb, 32'hc2b54d43, 32'hc10aa1c4, 32'h408d4708};
test_label[3277] = '{32'hc272daf1};
test_output[3277] = '{32'h42ed4a52};
/*############ DEBUG ############
test_input[26216:26223] = '{-93.7389520012, -32.286045943, -60.7138112386, 57.9313440562, -87.4507680854, -90.6509000061, -8.66449322713, 4.41492074697};
test_label[3277] = '{-60.7138112386};
test_output[3277] = '{118.645155295};
############ END DEBUG ############*/
test_input[26224:26231] = '{32'h42c1e9e3, 32'h42073fb4, 32'h4205f954, 32'hc2466a97, 32'hc270cb3b, 32'hc2945e2c, 32'h41a0e30e, 32'h4297fa27};
test_label[3278] = '{32'h4205f954};
test_output[3278] = '{32'h427dda71};
/*############ DEBUG ############
test_input[26224:26231] = '{96.9568075002, 33.8122118007, 33.493484135, -49.6040921609, -60.1984682613, -74.1839308404, 20.1108660894, 75.9885784814};
test_label[3278] = '{33.493484135};
test_output[3278] = '{63.463323366};
############ END DEBUG ############*/
test_input[26232:26239] = '{32'hc2bebd9d, 32'h4248d9ca, 32'h4208f24d, 32'h42030581, 32'hc2ba2a61, 32'h41c88e32, 32'h41c9f202, 32'h42b93063};
test_label[3279] = '{32'h4208f24d};
test_output[3279] = '{32'h42696e78};
/*############ DEBUG ############
test_input[26232:26239] = '{-95.3703395997, 50.2126851373, 34.2366231866, 32.7553760617, -93.0827733959, 25.069432025, 25.243167345, 92.5945034705};
test_label[3279] = '{34.2366231866};
test_output[3279] = '{58.3578802839};
############ END DEBUG ############*/
test_input[26240:26247] = '{32'h4272cb35, 32'h429ec46f, 32'hc2af90bb, 32'h3fea4001, 32'h422c3d84, 32'h41ad1b49, 32'h424a675d, 32'hc1abeb0f};
test_label[3280] = '{32'h3fea4001};
test_output[3280] = '{32'h429b1b6f};
/*############ DEBUG ############
test_input[26240:26247] = '{60.6984450838, 79.3836561286, -87.7826749903, 1.83007821697, 43.0600733179, 21.6383231494, 50.6009415416, -21.4897754292};
test_label[3280] = '{1.83007821697};
test_output[3280] = '{77.5535779193};
############ END DEBUG ############*/
test_input[26248:26255] = '{32'hc2163e47, 32'h42ac3c5b, 32'h424ea54c, 32'h425c51d3, 32'hc1cef567, 32'h427a4240, 32'h42567cc6, 32'h42b1f980};
test_label[3281] = '{32'hc2163e47};
test_output[3281] = '{32'h42fd34e5};
/*############ DEBUG ############
test_input[26248:26255] = '{-37.5608187667, 86.1178794724, 51.6614215444, 55.0799071426, -25.8698245919, 62.5646965674, 53.6218482153, 88.9873075105};
test_label[3281] = '{-37.5608187667};
test_output[3281] = '{126.603306804};
############ END DEBUG ############*/
test_input[26256:26263] = '{32'h422f7f43, 32'hc27053fa, 32'hc1de8ff5, 32'h41c08d5c, 32'h4293aaa1, 32'h427268b6, 32'hc2a91ad0, 32'h421897cf};
test_label[3282] = '{32'hc2a91ad0};
test_output[3282] = '{32'h431e62b8};
/*############ DEBUG ############
test_input[26256:26263] = '{43.8742774091, -60.0820075579, -27.8202916427, 24.0690222855, 73.8332573786, 60.602256877, -84.5523677393, 38.1482524422};
test_label[3282] = '{-84.5523677393};
test_output[3282] = '{158.385626912};
############ END DEBUG ############*/
test_input[26264:26271] = '{32'h42271dc7, 32'hbec306f3, 32'hc1ef633a, 32'h42605fcb, 32'hc2866350, 32'hc24a4ac1, 32'h420764bd, 32'hc0e89bc6};
test_label[3283] = '{32'hbec306f3};
test_output[3283] = '{32'h4261e5d9};
/*############ DEBUG ############
test_input[26264:26271] = '{41.7790782021, -0.380912404469, -29.9234503882, 56.0935483524, -67.1939720208, -50.5730021875, 33.8483767628, -7.26901537491};
test_label[3283] = '{-0.380912404469};
test_output[3283] = '{56.4744613642};
############ END DEBUG ############*/
test_input[26272:26279] = '{32'hc218b211, 32'hc29124d0, 32'h42b5ae1f, 32'h4233c2d5, 32'h422b0e5a, 32'hc28ca611, 32'h41b4dd5b, 32'hc2958c23};
test_label[3284] = '{32'h4233c2d5};
test_output[3284] = '{32'h42379968};
/*############ DEBUG ############
test_input[26272:26279] = '{-38.1738938364, -72.5718980342, 90.8400792403, 44.9402669081, 42.764014152, -70.3243449518, 22.6080834475, -74.7737073988};
test_label[3284] = '{44.9402669081};
test_output[3284] = '{45.8998123322};
############ END DEBUG ############*/
test_input[26280:26287] = '{32'h42bbc9c5, 32'hc28256e2, 32'h4290d4a4, 32'hc147f397, 32'hc2413359, 32'hc1f8db0c, 32'hc2891d9a, 32'h402dfd14};
test_label[3285] = '{32'hc28256e2};
test_output[3285] = '{32'h431f1053};
/*############ DEBUG ############
test_input[26280:26287] = '{93.8940781178, -65.1696937611, 72.4153158204, -12.4969697186, -48.3001452594, -31.1069569192, -68.557812635, 2.71857169127};
test_label[3285] = '{-65.1696937611};
test_output[3285] = '{159.063771879};
############ END DEBUG ############*/
test_input[26288:26295] = '{32'hc28c2666, 32'hc1e2a3bc, 32'hc2985617, 32'hc09fe93c, 32'hc29750db, 32'h424d03d7, 32'h4298c40a, 32'h428042d3};
test_label[3286] = '{32'hc1e2a3bc};
test_output[3286] = '{32'h42d16cfa};
/*############ DEBUG ############
test_input[26288:26295] = '{-70.0749944754, -28.3299492164, -76.1681450119, -4.99722109873, -75.6579191149, 51.2537480795, 76.3828902044, 64.1305161588};
test_label[3286] = '{-28.3299492164};
test_output[3286] = '{104.712844195};
############ END DEBUG ############*/
test_input[26296:26303] = '{32'hc15f8266, 32'h40ba4da3, 32'hc2484180, 32'hc28ae1dc, 32'hc17e23ac, 32'hc259826c, 32'hc2ab2733, 32'hc1e0eed6};
test_label[3287] = '{32'hc1e0eed6};
test_output[3287] = '{32'h4207c11f};
/*############ DEBUG ############
test_input[26296:26303] = '{-13.9693354606, 5.8219772073, -50.0639664223, -69.4411346067, -15.8837085492, -54.3773663347, -85.5765629815, -28.1166194171};
test_label[3287] = '{-28.1166194171};
test_output[3287] = '{33.9385966273};
############ END DEBUG ############*/
test_input[26304:26311] = '{32'hc2b88c0a, 32'h422d7d2b, 32'h42028aa5, 32'h42bee83f, 32'h4299e7f6, 32'hc24a4e6a, 32'h42256c25, 32'h425f449f};
test_label[3288] = '{32'h4299e7f6};
test_output[3288] = '{32'h41940122};
/*############ DEBUG ############
test_input[26304:26311] = '{-92.2735103363, 43.3722353832, 32.6353948926, 95.4536020187, 76.9530495282, -50.5765776823, 41.3556081178, 55.8170143604};
test_label[3288] = '{76.9530495282};
test_output[3288] = '{18.5005524997};
############ END DEBUG ############*/
test_input[26312:26319] = '{32'hc286bd7a, 32'hc28a3ef9, 32'h4214b6f3, 32'hc183e866, 32'hc2b313c0, 32'hc2ab2cdd, 32'h429f0f66, 32'hc1f2661f};
test_label[3289] = '{32'hc2ab2cdd};
test_output[3289] = '{32'h43251e21};
/*############ DEBUG ############
test_input[26312:26319] = '{-67.3700699745, -69.1229944526, 37.1786604989, -16.4884751648, -89.5385732469, -85.5876201956, 79.5300738253, -30.2998645721};
test_label[3289] = '{-85.5876201956};
test_output[3289] = '{165.117694021};
############ END DEBUG ############*/
test_input[26320:26327] = '{32'h4271e695, 32'h425cffaa, 32'hc2c540df, 32'hc279523f, 32'hc29c9af6, 32'hc1ccf768, 32'hc1405182, 32'h41c68e45};
test_label[3290] = '{32'h4271e695};
test_output[3290] = '{32'h3bafbe2d};
/*############ DEBUG ############
test_input[26320:26327] = '{60.4751762109, 55.2496733294, -98.6267031274, -62.3303201947, -78.3026552792, -25.6208034564, -12.0198992385, 24.8194678964};
test_label[3290] = '{60.4751762109};
test_output[3290] = '{0.00536324700107};
############ END DEBUG ############*/
test_input[26328:26335] = '{32'h404cebef, 32'hc2bd8a7d, 32'h423a5d44, 32'h41c80128, 32'h41eeabff, 32'hc25cc98a, 32'hc13dbad9, 32'h4177893d};
test_label[3291] = '{32'h423a5d44};
test_output[3291] = '{32'h3364806f};
/*############ DEBUG ############
test_input[26328:26335] = '{3.20190032672, -94.7704818217, 46.5910778065, 25.0005642385, 29.8339833614, -55.1968168966, -11.858116683, 15.4710058518};
test_label[3291] = '{46.5910778065};
test_output[3291] = '{5.32021968422e-08};
############ END DEBUG ############*/
test_input[26336:26343] = '{32'hc2811440, 32'h42c34a60, 32'hc2abb323, 32'hbff9fdae, 32'hc2c424b6, 32'h41b4abad, 32'hc2895d30, 32'h3f913a60};
test_label[3292] = '{32'hc2abb323};
test_output[3292] = '{32'h43377ec1};
/*############ DEBUG ############
test_input[26336:26343] = '{-64.5395488189, 97.6452610676, -85.8498778715, -1.95305413385, -98.0716999915, 22.5838260445, -68.6820104907, 1.13459401043};
test_label[3292] = '{-85.8498778715};
test_output[3292] = '{183.495138939};
############ END DEBUG ############*/
test_input[26344:26351] = '{32'hc2112598, 32'h42a3bc78, 32'h41ba4c7a, 32'hc2a70cd4, 32'h41f1462a, 32'hc2b99adb, 32'h41b00731, 32'h419fa260};
test_label[3293] = '{32'hc2112598};
test_output[3293] = '{32'h42ec4f44};
/*############ DEBUG ############
test_input[26344:26351] = '{-36.286712421, 81.8681035317, 23.2873420216, -83.5250579303, 30.1592596425, -92.802455796, 22.0035106345, 19.9542839706};
test_label[3293] = '{-36.286712421};
test_output[3293] = '{118.154815953};
############ END DEBUG ############*/
test_input[26352:26359] = '{32'hc144e39c, 32'hc2ada276, 32'hc2ba7acd, 32'hc24f5ddd, 32'h42a88315, 32'h42c04422, 32'h42989967, 32'hc11ee631};
test_label[3294] = '{32'hc144e39c};
test_output[3294] = '{32'h42d8e097};
/*############ DEBUG ############
test_input[26352:26359] = '{-12.3055688136, -86.8173078995, -93.239845912, -51.8416628304, 84.2560226973, 96.1330756958, 76.2996143456, -9.93119928399};
test_label[3294] = '{-12.3055688136};
test_output[3294] = '{108.43865146};
############ END DEBUG ############*/
test_input[26360:26367] = '{32'hc2a2e831, 32'hc192dfbb, 32'hc29db5f1, 32'hc243dc1b, 32'hc1acbdb8, 32'hc27993b3, 32'h4044385d, 32'hc127040e};
test_label[3295] = '{32'hc29db5f1};
test_output[3295] = '{32'h42a3d7b4};
/*############ DEBUG ############
test_input[26360:26367] = '{-81.4534971552, -18.3592437617, -78.8553565197, -48.9649476452, -21.5926353677, -62.3942373668, 3.0659401277, -10.4384895061};
test_label[3295] = '{-78.8553565197};
test_output[3295] = '{81.9212980128};
############ END DEBUG ############*/
test_input[26368:26375] = '{32'hc2b1f130, 32'hc29b0082, 32'hc1c7edbd, 32'h4283c360, 32'h42a37d90, 32'h42c2c244, 32'h42c66a4c, 32'h42c54578};
test_label[3296] = '{32'hc1c7edbd};
test_output[3296] = '{32'h42f97cee};
/*############ DEBUG ############
test_input[26368:26375] = '{-88.9710714028, -77.5009943191, -24.9910822066, 65.8815926725, 81.7452421785, 97.3794268009, 99.2076119973, 98.6356801767};
test_label[3296] = '{-24.9910822066};
test_output[3296] = '{124.744001817};
############ END DEBUG ############*/
test_input[26376:26383] = '{32'h41981283, 32'h4280fd8b, 32'h42965934, 32'hc1e37915, 32'hc29d96d8, 32'h4186f37b, 32'hc1a7b6cf, 32'hc2623cc4};
test_label[3297] = '{32'hc1e37915};
test_output[3297] = '{32'h42cf377c};
/*############ DEBUG ############
test_input[26376:26383] = '{19.0090394551, 64.4951975916, 75.1742230397, -28.4341211776, -78.7946149403, 16.8688876177, -20.9642624949, -56.5593401079};
test_label[3297] = '{-28.4341211776};
test_output[3297] = '{103.60836724};
############ END DEBUG ############*/
test_input[26384:26391] = '{32'h404b522e, 32'hc2b50be9, 32'hbc849db0, 32'h4220e1ca, 32'hc1a6e8a0, 32'hc2693d98, 32'hc270794f, 32'h42a66c7e};
test_label[3298] = '{32'hbc849db0};
test_output[3298] = '{32'h42a674c8};
/*############ DEBUG ############
test_input[26384:26391] = '{3.176890869, -90.5232629304, -0.0161884723089, 40.2204987708, -20.8635866584, -58.3101482935, -60.1184671739, 83.2118999413};
test_label[3298] = '{-0.0161884723089};
test_output[3298] = '{83.2280884136};
############ END DEBUG ############*/
test_input[26392:26399] = '{32'h420a520f, 32'h42bb0572, 32'hc205a4c1, 32'h426d8fe6, 32'h422bfe24, 32'hc0a64cd4, 32'hc215dd80, 32'h42a90223};
test_label[3299] = '{32'h426d8fe6};
test_output[3299] = '{32'h42087b1e};
/*############ DEBUG ############
test_input[26392:26399] = '{34.5801369101, 93.5106371818, -33.4108908129, 59.390527624, 42.9981844746, -5.19687843128, -37.4663076692, 84.5041767884};
test_label[3299] = '{59.390527624};
test_output[3299] = '{34.1202321654};
############ END DEBUG ############*/
test_input[26400:26407] = '{32'h429efd23, 32'h42693170, 32'hc1e35635, 32'hc237a72e, 32'hc20b7a02, 32'h42101dce, 32'h41466be9, 32'hc20e8dfa};
test_label[3300] = '{32'hc20b7a02};
test_output[3300] = '{32'h42e4ba24};
/*############ DEBUG ############
test_input[26400:26407] = '{79.4944053505, 58.2982790236, -28.4170925029, -45.9132631587, -34.8691486848, 36.0291065795, 12.4013457154, -35.6386483071};
test_label[3300] = '{-34.8691486848};
test_output[3300] = '{114.363554036};
############ END DEBUG ############*/
test_input[26408:26415] = '{32'hc141b37d, 32'h408d49cf, 32'h42449892, 32'h428ecb97, 32'hc249b0c7, 32'hc231f554, 32'hc2a1bf8c, 32'h41fcd1ee};
test_label[3301] = '{32'h41fcd1ee};
test_output[3301] = '{32'h421f2e37};
/*############ DEBUG ############
test_input[26408:26415] = '{-12.1063207027, 4.41525996876, 49.1489952927, 71.3976387053, -50.4226348646, -44.4895784685, -80.8741170653, 31.602505203};
test_label[3301] = '{31.602505203};
test_output[3301] = '{39.7951335025};
############ END DEBUG ############*/
test_input[26416:26423] = '{32'h4095be16, 32'hc2a95b68, 32'hc2afa6f6, 32'hc1a467aa, 32'hc23b0483, 32'h41de9450, 32'h42a34b55, 32'hc1faed03};
test_label[3302] = '{32'h41de9450};
test_output[3302] = '{32'h42574c82};
/*############ DEBUG ############
test_input[26416:26423] = '{4.67945366318, -84.67853085, -87.8260959207, -20.550617735, -46.7544046595, 27.8224179522, 81.6471315217, -31.365728244};
test_label[3302] = '{27.8224179522};
test_output[3302] = '{53.8247135695};
############ END DEBUG ############*/
test_input[26424:26431] = '{32'h42a006d4, 32'h42359021, 32'h4284b8c2, 32'hc0cce2d6, 32'h42a517d7, 32'hc287a194, 32'hc20a4094, 32'h40b88456};
test_label[3303] = '{32'hc0cce2d6};
test_output[3303] = '{32'h42b20d23};
/*############ DEBUG ############
test_input[26424:26431] = '{80.013339202, 45.3907498999, 66.360857509, -6.40269013544, 82.546560845, -67.8155837174, -34.5630640779, 5.76615426129};
test_label[3303] = '{-6.40269013544};
test_output[3303] = '{89.0256589926};
############ END DEBUG ############*/
test_input[26432:26439] = '{32'h42222e37, 32'hc0460f33, 32'h4280f605, 32'hc2208f32, 32'hc1258f40, 32'h4122db5d, 32'hc2a4f533, 32'h42bf11d2};
test_label[3304] = '{32'h4280f605};
test_output[3304] = '{32'h41f86f33};
/*############ DEBUG ############
test_input[26432:26439] = '{40.5451310604, -3.0946775888, 64.4805092508, -40.1398391847, -10.3474729474, 10.1785554288, -82.4789021464, 95.5348051193};
test_label[3304] = '{64.4805092508};
test_output[3304] = '{31.0542958686};
############ END DEBUG ############*/
test_input[26440:26447] = '{32'hc1e278cf, 32'hc287d235, 32'h426ebdd2, 32'h41dcd41e, 32'hc1221a4e, 32'hc25889aa, 32'h42a73b29, 32'h41f6f303};
test_label[3305] = '{32'h41f6f303};
test_output[3305] = '{32'h4252fcd1};
/*############ DEBUG ############
test_input[26440:26447] = '{-28.3089889574, -67.9105606596, 59.6853697579, 27.6035731872, -10.1314225153, -54.1344392049, 83.6155485807, 30.8686574864};
test_label[3305] = '{30.8686574864};
test_output[3305] = '{52.7468910943};
############ END DEBUG ############*/
test_input[26448:26455] = '{32'h42506d8b, 32'hc14ce4f1, 32'h4247b14f, 32'h428b42ad, 32'hc2858f0b, 32'h42c3d5ef, 32'hc1eba5ea, 32'hc1aa324c};
test_label[3306] = '{32'h428b42ad};
test_output[3306] = '{32'h41e24d05};
/*############ DEBUG ############
test_input[26448:26455] = '{52.1069771224, -12.8058934392, 49.9231530961, 69.6302271871, -66.7793837827, 97.9178352451, -29.4560122166, -21.2745589761};
test_label[3306] = '{69.6302271871};
test_output[3306] = '{28.287608058};
############ END DEBUG ############*/
test_input[26456:26463] = '{32'hc29f6399, 32'h428d6439, 32'hc2ac3c18, 32'hc2a812c8, 32'h420d00ac, 32'h425ec855, 32'h42bd9f09, 32'h42c3e7a6};
test_label[3307] = '{32'hc2a812c8};
test_output[3307] = '{32'h4336080b};
/*############ DEBUG ############
test_input[26456:26463] = '{-79.6945280371, 70.6957505009, -86.1173681856, -84.0366799949, 35.2506563959, 55.6956380742, 94.8106157321, 97.9524417327};
test_label[3307] = '{-84.0366799949};
test_output[3307] = '{182.031418316};
############ END DEBUG ############*/
test_input[26464:26471] = '{32'hc2bb89b0, 32'h428339f4, 32'hc2bdcc8e, 32'hc228f55c, 32'h4290e9e6, 32'h42934100, 32'h4237d8f0, 32'h41a8ee0e};
test_label[3308] = '{32'hc2bdcc8e};
test_output[3308] = '{32'h4328cc08};
/*############ DEBUG ############
test_input[26464:26471] = '{-93.7689208805, 65.6131915623, -94.8995187809, -42.2396079282, 72.4568338025, 73.6269534229, 45.9618540241, 21.1162372458};
test_label[3308] = '{-94.8995187809};
test_output[3308] = '{168.797003561};
############ END DEBUG ############*/
test_input[26472:26479] = '{32'hc1b62d49, 32'h4060345f, 32'hc19c67e7, 32'h4175b60c, 32'hc183a6ae, 32'h42b07b86, 32'hc20b530a, 32'h40beb10f};
test_label[3309] = '{32'hc20b530a};
test_output[3309] = '{32'h42f6250b};
/*############ DEBUG ############
test_input[26472:26479] = '{-22.7721118196, 3.50319648906, -19.550733289, 15.3569445745, -16.4563858189, 88.2412559753, -34.8310910468, 5.95911353944};
test_label[3309] = '{-34.8310910468};
test_output[3309] = '{123.072347022};
############ END DEBUG ############*/
test_input[26480:26487] = '{32'h42baa806, 32'h428466ac, 32'hc243686d, 32'h42bd3dad, 32'hc2766d42, 32'hc209069a, 32'h418b7f33, 32'hc240deb3};
test_label[3310] = '{32'h418b7f33};
test_output[3310] = '{32'h429ada1f};
/*############ DEBUG ############
test_input[26480:26487] = '{93.3281739444, 66.2005305248, -48.8519771423, 94.6204635841, -61.606697717, -34.256445604, 17.4371096601, -48.217478441};
test_label[3310] = '{17.4371096601};
test_output[3310] = '{77.4260186773};
############ END DEBUG ############*/
test_input[26488:26495] = '{32'hc2935b19, 32'h41924745, 32'hc2ac8cb8, 32'hc29b7de9, 32'h427c0783, 32'hc260866e, 32'h4291cdc3, 32'h41dba7ec};
test_label[3311] = '{32'hc2ac8cb8};
test_output[3311] = '{32'h431f2d41};
/*############ DEBUG ############
test_input[26488:26495] = '{-73.6779263097, 18.2847999604, -86.274842485, -77.7459178896, 63.0073362572, -56.1312775932, 72.901874705, 27.4569924375};
test_label[3311] = '{-86.274842485};
test_output[3311] = '{159.176767638};
############ END DEBUG ############*/
test_input[26496:26503] = '{32'hc28a974a, 32'hc23808be, 32'hc2881826, 32'hc25bc808, 32'h42130bd2, 32'hc084df8f, 32'h42228268, 32'h427068d7};
test_label[3312] = '{32'hc2881826};
test_output[3312] = '{32'h43002648};
/*############ DEBUG ############
test_input[26496:26503] = '{-69.2954882258, -46.0085387719, -68.0471620208, -54.9453441921, 36.7615436194, -4.15229005006, 40.6273497674, 60.1023816149};
test_label[3312] = '{-68.0471620208};
test_output[3312] = '{128.149543639};
############ END DEBUG ############*/
test_input[26504:26511] = '{32'h414b5044, 32'h42a244ce, 32'hc2670e08, 32'h4276c27b, 32'h424f6bd2, 32'h426f6b00, 32'h41af53c0, 32'hc225012d};
test_label[3313] = '{32'hc2670e08};
test_output[3313] = '{32'h430ae5e9};
/*############ DEBUG ############
test_input[26504:26511] = '{12.7070958774, 81.1343808761, -57.7637037521, 61.689923702, 51.8552915788, 59.8544904412, 21.9158933305, -41.2511487874};
test_label[3313] = '{-57.7637037521};
test_output[3313] = '{138.898084632};
############ END DEBUG ############*/
test_input[26512:26519] = '{32'h4212eef1, 32'h42597c61, 32'h41c8288b, 32'h429ff8af, 32'h41f71157, 32'h41e44f62, 32'h4280b6f7, 32'hc2c72628};
test_label[3314] = '{32'h41f71157};
test_output[3314] = '{32'h424468b2};
/*############ DEBUG ############
test_input[26512:26519] = '{36.7333408748, 54.3714653908, 25.0197963838, 79.985708857, 30.8834671977, 28.5387605636, 64.357352136, -99.5745233891};
test_label[3314] = '{30.8834671977};
test_output[3314] = '{49.1022418225};
############ END DEBUG ############*/
test_input[26520:26527] = '{32'h42c38e0b, 32'h429fbc5a, 32'h41ec1fb8, 32'hc1ef803b, 32'hc2a4149d, 32'h41d785fb, 32'hc2847256, 32'hc2235ee4};
test_label[3315] = '{32'hc2235ee4};
test_output[3315] = '{32'h430a9ebe};
/*############ DEBUG ############
test_input[26520:26527] = '{97.7774249457, 79.8678758106, 29.5154881046, -29.9376131374, -82.0402627566, 26.9404209822, -66.2233099096, -40.8426671331};
test_label[3315] = '{-40.8426671331};
test_output[3315] = '{138.620092095};
############ END DEBUG ############*/
test_input[26528:26535] = '{32'h426f0d0b, 32'hc2b35fae, 32'hc2a28601, 32'hc2115362, 32'h42a4e5e0, 32'h41db2bfc, 32'h4270da6e, 32'hc29fb493};
test_label[3316] = '{32'h41db2bfc};
test_output[3316] = '{32'h425c35c2};
/*############ DEBUG ############
test_input[26528:26535] = '{59.7627382192, -89.6868726356, -81.2617245081, -36.3314273872, 82.4489753885, 27.3964762844, 60.21330893, -79.8526818047};
test_label[3316] = '{27.3964762844};
test_output[3316] = '{55.0524991045};
############ END DEBUG ############*/
test_input[26536:26543] = '{32'hc1c12253, 32'hc099d01e, 32'h41d3e6ae, 32'h42566ca3, 32'h4286d750, 32'hc293869d, 32'h42b51dfe, 32'h4167dc01};
test_label[3317] = '{32'hc099d01e};
test_output[3317] = '{32'h42bebb00};
/*############ DEBUG ############
test_input[26536:26543] = '{-24.1417600814, -4.80665507752, 26.4876364534, 53.6060904536, 67.4205345081, -73.7629148586, 90.558582264, 14.4912122427};
test_label[3317] = '{-4.80665507752};
test_output[3317] = '{95.3652373416};
############ END DEBUG ############*/
test_input[26544:26551] = '{32'h429214e1, 32'h4183aaca, 32'hc096c9f5, 32'h42823be7, 32'h428ce5e2, 32'h429bd89a, 32'hc18d9483, 32'hc0053656};
test_label[3318] = '{32'h429214e1};
test_output[3318] = '{32'h409c7e19};
/*############ DEBUG ############
test_input[26544:26551] = '{73.040775483, 16.4583938919, -4.71215291198, 65.1169961917, 70.4489869028, 77.9230510836, -17.697515249, -2.0814413494};
test_label[3318] = '{73.040775483};
test_output[3318] = '{4.89039267457};
############ END DEBUG ############*/
test_input[26552:26559] = '{32'h42860efb, 32'hc27386bc, 32'hc15f01ca, 32'hc2b26602, 32'hc1c692e7, 32'hc253fbd7, 32'hc0fec6f9, 32'h428d5c5d};
test_label[3319] = '{32'hc253fbd7};
test_output[3319] = '{32'h42f76768};
/*############ DEBUG ############
test_input[26552:26559] = '{67.0292617381, -60.8815773515, -13.9379364146, -89.1992322459, -24.821730585, -52.9959385498, -7.96178858132, 70.680393844};
test_label[3319] = '{-52.9959385498};
test_output[3319] = '{123.701962831};
############ END DEBUG ############*/
test_input[26560:26567] = '{32'h427e6883, 32'h429ba9aa, 32'h408152ee, 32'hc1f183cb, 32'h42264f17, 32'hc1ce9a03, 32'h42ae41f1, 32'hc2bd7d03};
test_label[3320] = '{32'hc1f183cb};
test_output[3320] = '{32'h42eaa2f0};
/*############ DEBUG ############
test_input[26560:26567] = '{63.6020611081, 77.8313750456, 4.04137303356, -30.189351227, 41.5772355931, -25.8252012048, 87.1287911649, -94.7441639982};
test_label[3320] = '{-30.189351227};
test_output[3320] = '{117.318234048};
############ END DEBUG ############*/
test_input[26568:26575] = '{32'h42c2ce28, 32'hc2961567, 32'hc21d7dee, 32'h4177b22a, 32'h42c7f024, 32'h429d350e, 32'hc1c62c78, 32'h42b3adaf};
test_label[3321] = '{32'h4177b22a};
test_output[3321] = '{32'h42a91fc7};
/*############ DEBUG ############
test_input[26568:26575] = '{97.402645733, -75.0417993652, -39.3729772839, 15.4809972241, 99.9690211026, 78.603626006, -24.7717128069, 89.8392261008};
test_label[3321] = '{15.4809972241};
test_output[3321] = '{84.5620670892};
############ END DEBUG ############*/
test_input[26576:26583] = '{32'h42893489, 32'h42092d2d, 32'h42bff0ee, 32'hc2a50fe0, 32'h41d33ce3, 32'hc271ceaa, 32'hc2befce3, 32'hc2ac9eb0};
test_label[3322] = '{32'hc2a50fe0};
test_output[3322] = '{32'h43328067};
/*############ DEBUG ############
test_input[26576:26583] = '{68.602609094, 34.2941173353, 95.9705656102, -82.5310069041, 26.4047300477, -60.4518189278, -95.4939169758, -86.3099359065};
test_label[3322] = '{-82.5310069041};
test_output[3322] = '{178.501572514};
############ END DEBUG ############*/
test_input[26584:26591] = '{32'h42847fc7, 32'hc28c0bed, 32'h427f3205, 32'h4019b2e6, 32'hc0835712, 32'h427e2e66, 32'hc14188a3, 32'hc0d0d60b};
test_label[3323] = '{32'h4019b2e6};
test_output[3323] = '{32'h427ff64b};
/*############ DEBUG ############
test_input[26584:26591] = '{66.2495669407, -70.0232933306, 63.7988473984, 2.40154411431, -4.10437893697, 63.5453127336, -12.0958588416, -6.5261281203};
test_label[3323] = '{2.40154411431};
test_output[3323] = '{63.9905216555};
############ END DEBUG ############*/
test_input[26592:26599] = '{32'h42c4036a, 32'h41933054, 32'hc29072d5, 32'h42242e1d, 32'h413cd2ac, 32'hc2beab3a, 32'h428eab34, 32'h42a3d238};
test_label[3324] = '{32'hc2beab3a};
test_output[3324] = '{32'h43415752};
/*############ DEBUG ############
test_input[26592:26599] = '{98.0066644643, 18.3985974419, -72.2242785897, 41.0450342211, 11.8014334245, -95.3344249889, 71.3343792566, 81.9105802606};
test_label[3324] = '{-95.3344249889};
test_output[3324] = '{193.341089555};
############ END DEBUG ############*/
test_input[26600:26607] = '{32'hc291ec8c, 32'h428ae7bf, 32'hc29a29a0, 32'hc1e713b6, 32'hc285546a, 32'hbed04190, 32'hc23a4277, 32'h423a9871};
test_label[3325] = '{32'hbed04190};
test_output[3325] = '{32'h428bb801};
/*############ DEBUG ############
test_input[26600:26607] = '{-72.9620079892, 69.4526326226, -77.0812988087, -28.8846253361, -66.6648702731, -0.406750198782, -46.5649074774, 46.6488687702};
test_label[3325] = '{-0.406750198782};
test_output[3325] = '{69.8593828215};
############ END DEBUG ############*/
test_input[26608:26615] = '{32'hc20a419e, 32'hc1d8785e, 32'hc2b07f4b, 32'h421ff468, 32'h426e999f, 32'hc2a48c2d, 32'hc29f9aca, 32'h425acf0d};
test_label[3326] = '{32'h421ff468};
test_output[3326] = '{32'h419d58eb};
/*############ DEBUG ############
test_input[26608:26615] = '{-34.5640782822, -27.0587739303, -88.2486164117, 39.9886770563, 59.650020522, -82.2737792155, -79.8023224187, 54.7021988052};
test_label[3326] = '{39.9886770563};
test_output[3326] = '{19.6684172456};
############ END DEBUG ############*/
test_input[26616:26623] = '{32'hc2174265, 32'h42598bf4, 32'hc28ac281, 32'h423f13eb, 32'hc2c4b747, 32'hc20f15ca, 32'hc2b02564, 32'h425a16de};
test_label[3327] = '{32'hc2b02564};
test_output[3327] = '{32'h430f393e};
/*############ DEBUG ############
test_input[26616:26623] = '{-37.8148385636, 54.3866725956, -69.3798873827, 47.7694523778, -98.3579619457, -35.7712766159, -88.0730318204, 54.5223325008};
test_label[3327] = '{-88.0730318204};
test_output[3327] = '{143.223603336};
############ END DEBUG ############*/
test_input[26624:26631] = '{32'h42c6336d, 32'hc28e5ce2, 32'h42a4fde8, 32'h41967809, 32'h417df776, 32'h427445ce, 32'hc13f2c3b, 32'hc295a9e2};
test_label[3328] = '{32'h42c6336d};
test_output[3328] = '{32'h338407cc};
/*############ DEBUG ############
test_input[26624:26631] = '{99.1004402584, -71.1814085838, 82.4959102693, 18.8086116351, 15.8729151834, 61.068166955, -11.948298721, -74.8318043058};
test_label[3328] = '{99.1004402584};
test_output[3328] = '{6.14814692516e-08};
############ END DEBUG ############*/
test_input[26632:26639] = '{32'h4203c837, 32'hc1c363f3, 32'hbfa789f8, 32'h41b049ae, 32'h429f1ecc, 32'h42bb0bb6, 32'hbd8ceaf0, 32'hc2045c29};
test_label[3329] = '{32'hbfa789f8};
test_output[3329] = '{32'h42bda9de};
/*############ DEBUG ############
test_input[26632:26639] = '{32.9455241121, -24.4238027658, -1.30889796952, 22.0359767337, 79.560152091, 93.5228761829, -0.0688074832539, -33.0899990152};
test_label[3329] = '{-1.30889796952};
test_output[3329] = '{94.8317750155};
############ END DEBUG ############*/
test_input[26640:26647] = '{32'h42ad1a04, 32'h42af8ba3, 32'h422a3508, 32'h411d2620, 32'h41962138, 32'hc238cb21, 32'hc27845ff, 32'h429e97f8};
test_label[3330] = '{32'hc238cb21};
test_output[3330] = '{32'h43063ac1};
/*############ DEBUG ############
test_input[26640:26647] = '{86.5508103648, 87.7727273772, 42.5517875977, 9.82180742536, 18.7662192147, -46.1983693382, -62.0683566519, 79.2968163703};
test_label[3330] = '{-46.1983693382};
test_output[3330] = '{134.229509474};
############ END DEBUG ############*/
test_input[26648:26655] = '{32'h425322ce, 32'h42836e87, 32'h423642f7, 32'h42b40e47, 32'hc2314180, 32'h423f2984, 32'h427d3872, 32'h42791693};
test_label[3331] = '{32'h423f2984};
test_output[3331] = '{32'h4228f30b};
/*############ DEBUG ############
test_input[26648:26655] = '{52.7839876917, 65.7158762265, 45.5653935159, 90.0278861796, -44.3139637654, 47.7905407509, 63.305122749, 62.2720469214};
test_label[3331] = '{47.7905407509};
test_output[3331] = '{42.2373454287};
############ END DEBUG ############*/
test_input[26656:26663] = '{32'hc28cb7cb, 32'hc254df1d, 32'hc2193d44, 32'h420032f2, 32'h41ca1c03, 32'hc117ef9f, 32'hc2b42cc7, 32'h42067746};
test_label[3332] = '{32'hc117ef9f};
test_output[3332] = '{32'h422d357f};
/*############ DEBUG ############
test_input[26656:26663] = '{-70.3589727281, -53.2178830447, -38.3098294436, 32.0497495786, 25.2636776293, -9.4960012738, -90.0874570073, 33.6164779553};
test_label[3332] = '{-9.4960012738};
test_output[3332] = '{43.30224193};
############ END DEBUG ############*/
test_input[26664:26671] = '{32'hc27cc83f, 32'h426be7cf, 32'h41792ee9, 32'hc1c5e5b1, 32'h42c42dbc, 32'h42a3eef2, 32'hc2a6921b, 32'h41f00f5d};
test_label[3333] = '{32'hc27cc83f};
test_output[3333] = '{32'h432148ee};
/*############ DEBUG ############
test_input[26664:26671] = '{-63.195551405, 58.976375513, 15.5739524003, -24.7371543364, 98.0893241201, 81.9666933431, -83.2853628061, 30.0075007318};
test_label[3333] = '{-63.195551405};
test_output[3333] = '{161.284875625};
############ END DEBUG ############*/
test_input[26672:26679] = '{32'hbf146db1, 32'hc26fcf70, 32'h41c2fe58, 32'h42380d64, 32'h41d7f2f0, 32'h42836f40, 32'h429e5713, 32'h42c14b0e};
test_label[3334] = '{32'h42836f40};
test_output[3334] = '{32'h41f76f37};
/*############ DEBUG ############
test_input[26672:26679] = '{-0.57979877114, -59.9525749128, 24.3741912947, 46.0130752289, 26.9936226589, 65.7172887829, 79.1700663044, 96.6465932274};
test_label[3334] = '{65.7172887829};
test_output[3334] = '{30.9293044702};
############ END DEBUG ############*/
test_input[26680:26687] = '{32'h423bc337, 32'h427da513, 32'h42029df7, 32'h41bad789, 32'h41b7d7c1, 32'h418fc184, 32'h428372ff, 32'h429c7661};
test_label[3335] = '{32'h423bc337};
test_output[3335] = '{32'h41fa5316};
/*############ DEBUG ############
test_input[26680:26687] = '{46.9406413223, 63.4112065866, 32.6542618724, 23.3552425343, 22.9803489465, 17.9694905703, 65.7245993236, 78.2312059304};
test_label[3335] = '{46.9406413223};
test_output[3335] = '{31.2905686764};
############ END DEBUG ############*/
test_input[26688:26695] = '{32'hc2010021, 32'hc1e9023b, 32'hc1acdf8e, 32'h42b8f49b, 32'hc2a3f7f5, 32'h425e76a2, 32'h4210ae3e, 32'hc2659e37};
test_label[3336] = '{32'h4210ae3e};
test_output[3336] = '{32'h42613af9};
/*############ DEBUG ############
test_input[26688:26695] = '{-32.2501259081, -29.1260884442, -21.6091583693, 92.4777468284, -81.984288134, 55.6158527056, 36.1701574965, -57.404506935};
test_label[3336] = '{36.1701574965};
test_output[3336] = '{56.3075893319};
############ END DEBUG ############*/
test_input[26696:26703] = '{32'h42286820, 32'hc16e6063, 32'h42b9e8cb, 32'h41d38aaf, 32'hc216ff5d, 32'hc21ee390, 32'h41db79cc, 32'h4176d224};
test_label[3337] = '{32'h41d38aaf};
test_output[3337] = '{32'h4285061f};
/*############ DEBUG ############
test_input[26696:26703] = '{42.1016857945, -14.8985319206, 92.954671307, 26.4427156549, -37.7493789478, -39.722229762, 27.434471789, 15.4263041978};
test_label[3337] = '{26.4427156549};
test_output[3337] = '{66.5119556522};
############ END DEBUG ############*/
test_input[26704:26711] = '{32'h426a452a, 32'h41f33921, 32'h42b1a77b, 32'hc28d2b1c, 32'h42a0e6a6, 32'h41ee4350, 32'h42bb6f5e, 32'hc2462f7c};
test_label[3338] = '{32'hc2462f7c};
test_output[3338] = '{32'h430f4579};
/*############ DEBUG ############
test_input[26704:26711] = '{58.5675448063, 30.4028943292, 88.8271129853, -70.5841987869, 80.450483069, 29.7828674533, 93.717512893, -49.5463733136};
test_label[3338] = '{-49.5463733136};
test_output[3338] = '{143.271378217};
############ END DEBUG ############*/
test_input[26712:26719] = '{32'h4206bc2b, 32'hc2a269ce, 32'hc0228479, 32'h41f9b31c, 32'h41e5e0e4, 32'h42a69f82, 32'hc234cd3c, 32'h42407c87};
test_label[3339] = '{32'h41f9b31c};
test_output[3339] = '{32'h42506575};
/*############ DEBUG ############
test_input[26712:26719] = '{33.6837592492, -81.2066525015, -2.53933554, 31.2124559297, 28.7348104154, 83.3115367418, -45.2004230165, 48.1216076735};
test_label[3339] = '{31.2124559297};
test_output[3339] = '{52.0990808121};
############ END DEBUG ############*/
test_input[26720:26727] = '{32'h42bef761, 32'hc2b597c0, 32'hc21ae79a, 32'h42285586, 32'hc22fc08a, 32'hc2170d26, 32'hc21b4749, 32'hc2b2085a};
test_label[3340] = '{32'h42bef761};
test_output[3340] = '{32'h80000000};
/*############ DEBUG ############
test_input[26720:26727] = '{95.4831605638, -90.7963868153, -38.726172713, 42.0835207087, -43.938026949, -37.7628386527, -38.8196157702, -89.0163091513};
test_label[3340] = '{95.4831605638};
test_output[3340] = '{-0.0};
############ END DEBUG ############*/
test_input[26728:26735] = '{32'hc2bc7a06, 32'hc288d095, 32'h429f4d2b, 32'h40a985a0, 32'hc2664c6e, 32'hc16afb0a, 32'hc256fc35, 32'h427af347};
test_label[3341] = '{32'hc2664c6e};
test_output[3341] = '{32'h430939b1};
/*############ DEBUG ############
test_input[26728:26735] = '{-94.2383305999, -68.4073849497, 79.6507212444, 5.29756157246, -57.5746371187, -14.6862885858, -53.7462958344, 62.7375754884};
test_label[3341] = '{-57.5746371187};
test_output[3341] = '{137.225358408};
############ END DEBUG ############*/
test_input[26736:26743] = '{32'h4229b9c5, 32'hc223acd0, 32'h42bbfa8c, 32'h42a6c890, 32'hc2a41493, 32'h42a97bf2, 32'hc2411d39, 32'hc221510a};
test_label[3342] = '{32'hc2a41493};
test_output[3342] = '{32'h43300797};
/*############ DEBUG ############
test_input[26736:26743] = '{42.4314139846, -40.9187628707, 93.9893497304, 83.3917202506, -82.0401810635, 84.7420814122, -48.278536712, -40.329139474};
test_label[3342] = '{-82.0401810635};
test_output[3342] = '{176.029652136};
############ END DEBUG ############*/
test_input[26744:26751] = '{32'h4289b2d9, 32'h4278ea4b, 32'h4241b729, 32'hc0510579, 32'h4273801a, 32'hc29de577, 32'hc2b8592d, 32'h42b49b8b};
test_label[3343] = '{32'hc29de577};
test_output[3343] = '{32'h43294081};
/*############ DEBUG ############
test_input[26744:26751] = '{68.849309969, 62.2288025224, 48.4288658341, -3.26595903454, 60.8750991101, -78.9481756527, -92.1741685684, 90.3037978588};
test_label[3343] = '{-78.9481756527};
test_output[3343] = '{169.251973512};
############ END DEBUG ############*/
test_input[26752:26759] = '{32'h425ed46b, 32'h426b213a, 32'hc1fd65f0, 32'h42b7df79, 32'h428328ec, 32'hc1efa4bf, 32'h4298659e, 32'h415e4a36};
test_label[3344] = '{32'h42b7df79};
test_output[3344] = '{32'h341d07bf};
/*############ DEBUG ############
test_input[26752:26759] = '{55.7074390752, 58.7824475768, -31.6747748056, 91.9364697325, 65.5799259871, -29.9554427199, 76.1984683853, 13.8931175412};
test_label[3344] = '{91.9364697325};
test_output[3344] = '{1.46245819712e-07};
############ END DEBUG ############*/
test_input[26760:26767] = '{32'hc24e6f62, 32'hc13a391f, 32'h42541ab6, 32'h42995560, 32'hbff6d495, 32'h409a6842, 32'h429de3b3, 32'hc01c7fde};
test_label[3345] = '{32'h409a6842};
test_output[3345] = '{32'h42946f24};
/*############ DEBUG ############
test_input[26760:26767] = '{-51.6087720493, -11.6389453832, 53.0260846269, 76.6667462984, -1.92836243592, 4.82522692479, 78.9447222876, -2.44530451161};
test_label[3345] = '{4.82522692479};
test_output[3345] = '{74.2170679276};
############ END DEBUG ############*/
test_input[26768:26775] = '{32'h425dc7ca, 32'hc2c2dd7a, 32'h429fb085, 32'h42551103, 32'hc1d87dcd, 32'hc23c55e2, 32'hc1a175d3, 32'h413ffd31};
test_label[3346] = '{32'h413ffd31};
test_output[3346] = '{32'h4287b0df};
/*############ DEBUG ############
test_input[26768:26775] = '{55.4451063943, -97.432572517, 79.84476806, 53.2666113833, -27.0614257458, -47.0838707978, -20.1825322717, 11.9993143482};
test_label[3346] = '{11.9993143482};
test_output[3346] = '{67.8454537119};
############ END DEBUG ############*/
test_input[26776:26783] = '{32'hc2bb3afc, 32'hc2b8d41b, 32'h41da59a2, 32'h42ab42e0, 32'hc2c75ad0, 32'h42a12721, 32'hc17c1e11, 32'hc2afa6d5};
test_label[3347] = '{32'h42a12721};
test_output[3347] = '{32'h40a1f006};
/*############ DEBUG ############
test_input[26776:26783] = '{-93.6152024282, -92.4142718636, 27.2937653595, 85.6306130711, -99.6773687384, 80.5764258082, -15.75734018, -87.825847176};
test_label[3347] = '{80.5764258082};
test_output[3347] = '{5.0605495327};
############ END DEBUG ############*/
test_input[26784:26791] = '{32'h412d7a57, 32'h40c69ed9, 32'h41911ce5, 32'hc21b1386, 32'hc2c7e318, 32'h42ae1c54, 32'h42aa5b4d, 32'hc2bc8b56};
test_label[3348] = '{32'h42aa5b4d};
test_output[3348] = '{32'h40013e16};
/*############ DEBUG ############
test_input[26784:26791] = '{10.8423680048, 6.20689066846, 18.1391093835, -38.7690675875, -99.943538766, 87.055327698, 85.178321765, -94.2721400367};
test_label[3348] = '{85.178321765};
test_output[3348] = '{2.01941450505};
############ END DEBUG ############*/
test_input[26792:26799] = '{32'hc299b59c, 32'h4196c6e8, 32'h42265179, 32'hc1692868, 32'hc278ed70, 32'hc2636712, 32'hc1bfb9bf, 32'h41d65165};
test_label[3349] = '{32'h4196c6e8};
test_output[3349] = '{32'h41b5dc09};
/*############ DEBUG ############
test_input[26792:26799] = '{-76.8547027088, 18.8471226558, 41.5795620633, -14.5723648389, -62.2318722067, -56.8506535245, -23.9656972527, 26.7897441473};
test_label[3349] = '{18.8471226558};
test_output[3349] = '{22.7324397851};
############ END DEBUG ############*/
test_input[26800:26807] = '{32'hc2429df2, 32'hc1c3e11b, 32'h41acd1b9, 32'h4240234e, 32'h429b21a3, 32'hc2b9fd5a, 32'hc1dcd4d0, 32'h409f5e3a};
test_label[3350] = '{32'hc2429df2};
test_output[3350] = '{32'h42fc709c};
/*############ DEBUG ############
test_input[26800:26807] = '{-48.6542439592, -24.4849141577, 21.6024027465, 48.0344765347, 77.5656996005, -92.9948307744, -27.6039129988, 4.98025239063};
test_label[3350] = '{-48.6542439592};
test_output[3350] = '{126.21994356};
############ END DEBUG ############*/
test_input[26808:26815] = '{32'hc23e06fb, 32'h424248c3, 32'hc1f9e0db, 32'hc2893581, 32'h412f9f3f, 32'h4272973b, 32'h42b0b564, 32'h41bf683a};
test_label[3351] = '{32'h42b0b564};
test_output[3351] = '{32'h2b828000};
/*############ DEBUG ############
test_input[26808:26815] = '{-47.5068157942, 48.5710551679, -31.2347930945, -68.6045032119, 10.9763780597, 60.6476877017, 88.354276254, 23.9258922536};
test_label[3351] = '{88.354276254};
test_output[3351] = '{9.27258270167e-13};
############ END DEBUG ############*/
test_input[26816:26823] = '{32'hc2c7747d, 32'h42a34283, 32'h422df92c, 32'hc2c6d1d7, 32'hc22dbf42, 32'h423b9d2a, 32'hc1a09a48, 32'h42a20678};
test_label[3352] = '{32'h422df92c};
test_output[3352] = '{32'h421a459b};
/*############ DEBUG ############
test_input[26816:26823] = '{-99.7275126868, 81.6299037162, 43.4933333526, -99.4098471938, -43.4367765811, 46.9034796741, -20.0753330138, 81.0126368477};
test_label[3352] = '{43.4933333526};
test_output[3352] = '{38.567973956};
############ END DEBUG ############*/
test_input[26824:26831] = '{32'hc18abd2e, 32'hc2107211, 32'hc21bbf0a, 32'hc2bede35, 32'h40c717b3, 32'hc16f3012, 32'hc288e021, 32'hc2afe2e5};
test_label[3353] = '{32'hc288e021};
test_output[3353] = '{32'h4295519c};
/*############ DEBUG ############
test_input[26824:26831] = '{-17.3423736006, -36.1113929155, -38.9365617447, -95.4339994427, 6.22164302797, -14.9492358211, -68.4377499174, -87.9431544298};
test_label[3353] = '{-68.4377499174};
test_output[3353] = '{74.6593929461};
############ END DEBUG ############*/
test_input[26832:26839] = '{32'hc284cb28, 32'h4238c924, 32'hc2a67dfd, 32'hc23cb7bc, 32'h3f479c52, 32'hc1c797bd, 32'hc22d46eb, 32'h416f9fb5};
test_label[3354] = '{32'hc284cb28};
test_output[3354] = '{32'h42e12fbb};
/*############ DEBUG ############
test_input[26832:26839] = '{-66.3967928323, 46.1964277627, -83.2460694341, -47.1794283063, 0.779729010062, -24.9490904039, -43.3192562831, 14.9764905458};
test_label[3354] = '{-66.3967928323};
test_output[3354] = '{112.593220595};
############ END DEBUG ############*/
test_input[26840:26847] = '{32'h42b53fab, 32'hc24a9bd2, 32'hc2a39dfb, 32'hc1ef24b7, 32'h418b4f87, 32'h425cdb15, 32'hc1d318c1, 32'hc16d197c};
test_label[3355] = '{32'hc24a9bd2};
test_output[3355] = '{32'h430d46ca};
/*############ DEBUG ############
test_input[26840:26847] = '{90.6243520478, -50.6521688229, -81.8085555069, -29.8929262259, 17.4138324905, 55.213949158, -26.387087448, -14.8187215925};
test_label[3355] = '{-50.6521688229};
test_output[3355] = '{141.276520871};
############ END DEBUG ############*/
test_input[26848:26855] = '{32'hc2938b66, 32'h4149ad43, 32'hc0bf4f84, 32'h4252b24e, 32'hc2b89ce5, 32'h4261931b, 32'h42a7a396, 32'hc2ac3610};
test_label[3356] = '{32'hc0bf4f84};
test_output[3356] = '{32'h42b3988f};
/*############ DEBUG ############
test_input[26848:26855] = '{-73.7722628753, 12.6048000739, -5.97845659547, 52.6741255119, -92.3064375884, 56.3936591309, 83.8195071569, -86.1055919271};
test_label[3356] = '{-5.97845659547};
test_output[3356] = '{89.7979637524};
############ END DEBUG ############*/
test_input[26856:26863] = '{32'hc14a0cff, 32'hc09b1cb5, 32'h4127e43a, 32'hc258d9b1, 32'hc28c0e5b, 32'h42aa3066, 32'hc29bcba5, 32'hc28521e7};
test_label[3357] = '{32'hc14a0cff};
test_output[3357] = '{32'h42c37206};
/*############ DEBUG ############
test_input[26856:26863] = '{-12.6281729176, -4.84725406925, 10.4932193211, -54.2125888276, -70.0280409344, 85.0945308346, -77.8977404724, -66.5662119334};
test_label[3357] = '{-12.6281729176};
test_output[3357] = '{97.7227037522};
############ END DEBUG ############*/
test_input[26864:26871] = '{32'hc10b5166, 32'h41cf98af, 32'h420b2409, 32'hc0c870ec, 32'hc2801747, 32'h41ef5ddb, 32'h41f6965a, 32'h42c5c104};
test_label[3358] = '{32'h420b2409};
test_output[3358] = '{32'h42802f00};
/*############ DEBUG ############
test_input[26864:26871] = '{-8.70737308767, 25.9495528537, 34.7851915145, -6.26378447871, -64.0454628094, 29.9208272343, 30.8234137697, 98.876985112};
test_label[3358] = '{34.7851915145};
test_output[3358] = '{64.0917935975};
############ END DEBUG ############*/
test_input[26872:26879] = '{32'h4119333d, 32'hc28148fb, 32'h42a37768, 32'h410da685, 32'h41f8e5a9, 32'h423cbe98, 32'h41b3bc92, 32'h40453a85};
test_label[3359] = '{32'h41f8e5a9};
test_output[3359] = '{32'h424a7bfb};
/*############ DEBUG ############
test_input[26872:26879] = '{9.57500966384, -64.6425385708, 81.733212345, 8.85315414381, 31.1121381242, 47.1861263487, 22.4670758636, 3.0816967592};
test_label[3359] = '{31.1121381242};
test_output[3359] = '{50.6210742209};
############ END DEBUG ############*/
test_input[26880:26887] = '{32'hc1f5840f, 32'hc236e921, 32'hc20a9c77, 32'hc20b85a7, 32'hc28a2a66, 32'hc2b1cd47, 32'h42b8fd14, 32'h4296877a};
test_label[3360] = '{32'h4296877a};
test_output[3360] = '{32'h4189d669};
/*############ DEBUG ############
test_input[26880:26887] = '{-30.6894813415, -45.7276663396, -34.6527988613, -34.8805214866, -69.082808361, -88.9009325267, 92.4942959062, 75.2646027729};
test_label[3360] = '{75.2646027729};
test_output[3360] = '{17.2296931662};
############ END DEBUG ############*/
test_input[26888:26895] = '{32'hc1d75d2e, 32'h421c2f07, 32'h41f60208, 32'hc2912580, 32'h428bef0a, 32'h41d78607, 32'hc138be72, 32'h42a71dd8};
test_label[3361] = '{32'h428bef0a};
test_output[3361] = '{32'h4159766f};
/*############ DEBUG ############
test_input[26888:26895] = '{-26.9204980291, 39.0459265267, 30.7509923929, -72.5732435832, 69.9668719261, 26.9404430737, -11.5464958556, 83.558284911};
test_label[3361] = '{69.9668719261};
test_output[3361] = '{13.5914142361};
############ END DEBUG ############*/
test_input[26896:26903] = '{32'hc127ce36, 32'hc2a0a9c0, 32'hc1253c9b, 32'hc2bb8355, 32'h41e3a916, 32'h41e66c6b, 32'h41283b92, 32'hc2abe15b};
test_label[3362] = '{32'hc2bb8355};
test_output[3362] = '{32'h42f63082};
/*############ DEBUG ############
test_input[26896:26903] = '{-10.4878445733, -80.3315418739, -10.3272966303, -93.7565090667, 28.4575623502, 28.8029383733, 10.5145431641, -85.9401456588};
test_label[3362] = '{-93.7565090667};
test_output[3362] = '{123.094743666};
############ END DEBUG ############*/
test_input[26904:26911] = '{32'h423412df, 32'hc231be10, 32'h427fef56, 32'hc2c63706, 32'h4273bb99, 32'hc25b4af1, 32'hc1aa50af, 32'h429ebf0e};
test_label[3363] = '{32'hc1aa50af};
test_output[3363] = '{32'h42c95339};
/*############ DEBUG ############
test_input[26904:26911] = '{45.0184269432, -44.4356072519, 63.9837267383, -99.1074676113, 60.9332009235, -54.8231855927, -21.2893959264, 79.3731509423};
test_label[3363] = '{-21.2893959264};
test_output[3363] = '{100.662547086};
############ END DEBUG ############*/
test_input[26912:26919] = '{32'hc2433640, 32'h423f7ecd, 32'h420fa60b, 32'h41016ae9, 32'hc2902022, 32'hc20239e3, 32'hc27ee304, 32'hc205064b};
test_label[3364] = '{32'h41016ae9};
test_output[3364] = '{32'h421f2415};
/*############ DEBUG ############
test_input[26912:26919] = '{-48.8029796762, 47.8738301011, 35.9121506277, 8.08860135614, -72.0627556003, -32.5565295257, -63.7216945786, -33.2561471591};
test_label[3364] = '{8.08860135614};
test_output[3364] = '{39.7852351292};
############ END DEBUG ############*/
test_input[26920:26927] = '{32'h41ae8d36, 32'hc2526c52, 32'hc21082c5, 32'hc2846ee7, 32'hc1754a6f, 32'hc276f1c4, 32'h415094db, 32'h425806a7};
test_label[3365] = '{32'hc2526c52};
test_output[3365] = '{32'h42d5397c};
/*############ DEBUG ############
test_input[26920:26927] = '{21.8189499956, -52.6057809224, -36.1277034828, -66.2166096056, -15.3306722374, -61.7360986444, 13.0363417809, 54.0064953186};
test_label[3365] = '{-52.6057809224};
test_output[3365] = '{106.612276241};
############ END DEBUG ############*/
test_input[26928:26935] = '{32'hc240df93, 32'h414bd666, 32'hc2841e5d, 32'h42960bca, 32'h428c9895, 32'h42b86065, 32'h41fe284a, 32'h3fbb05c6};
test_label[3366] = '{32'h42960bca};
test_output[3366] = '{32'h4189526d};
/*############ DEBUG ############
test_input[26928:26935] = '{-48.2183358065, 12.7398429324, -66.0593029283, 75.0230255592, 70.2980087732, 92.1882725899, 31.769673052, 1.46111365591};
test_label[3366] = '{75.0230255592};
test_output[3366] = '{17.1652470661};
############ END DEBUG ############*/
test_input[26936:26943] = '{32'h42c4284f, 32'h42348485, 32'hc2be0a91, 32'h422c68ae, 32'hc2c5b0cd, 32'hc044c2cc, 32'hc189a89d, 32'hc2947ef5};
test_label[3367] = '{32'hc044c2cc};
test_output[3367] = '{32'h42ca4e65};
/*############ DEBUG ############
test_input[26936:26943] = '{98.0787283177, 45.1294119091, -95.0206361947, 43.1022252866, -98.8453111513, -3.07438947526, -17.207330989, -74.2479640989};
test_label[3367] = '{-3.07438947526};
test_output[3367] = '{101.153117793};
############ END DEBUG ############*/
test_input[26944:26951] = '{32'h427a968e, 32'h41cd0309, 32'h426acd85, 32'hc1ceb6bb, 32'hc2bf124c, 32'hc1e19e8f, 32'h425d4efa, 32'hc248a31c};
test_label[3368] = '{32'h427a968e};
test_output[3368] = '{32'h3ca22024};
/*############ DEBUG ############
test_input[26944:26951] = '{62.6470274696, 25.6264814485, 58.7007040884, -25.8392231426, -95.535738067, -28.2024214976, 55.3271257371, -50.1592853031};
test_label[3368] = '{62.6470274696};
test_output[3368] = '{0.0197907169851};
############ END DEBUG ############*/
test_input[26952:26959] = '{32'h428ea825, 32'h427b58a9, 32'hc15a340c, 32'hc2c6cf3c, 32'h41ed0a7e, 32'h4288f939, 32'hc21a4d1d, 32'h422de4b9};
test_label[3369] = '{32'hc21a4d1d};
test_output[3369] = '{32'h42dbebd3};
/*############ DEBUG ############
test_input[26952:26959] = '{71.3284037492, 62.8365826325, -13.6377066732, -99.4047529822, 29.6301223105, 68.4867601708, -38.5753048994, 43.4733607463};
test_label[3369] = '{-38.5753048994};
test_output[3369] = '{109.96059439};
############ END DEBUG ############*/
test_input[26960:26967] = '{32'h42b6aa33, 32'h42b45b40, 32'h42be0c64, 32'h411515d2, 32'hc291f434, 32'hc28f0eff, 32'h41c49d82, 32'h40c53677};
test_label[3370] = '{32'h42b45b40};
test_output[3370] = '{32'h409c1a84};
/*############ DEBUG ############
test_input[26960:26967] = '{91.3324231837, 90.1782228128, 95.0241978964, 9.31782736754, -72.9769606449, -71.5292889966, 24.5769082495, 6.16289856442};
test_label[3370] = '{90.1782228128};
test_output[3370] = '{4.8782367084};
############ END DEBUG ############*/
test_input[26968:26975] = '{32'hc03e482d, 32'h42781127, 32'h429a8568, 32'h409d2d44, 32'h42c153e8, 32'h42c16bce, 32'h42ad8bfa, 32'h42462151};
test_label[3371] = '{32'h42ad8bfa};
test_output[3371] = '{32'h4129b761};
/*############ DEBUG ############
test_input[26968:26975] = '{-2.9731552829, 62.0167492282, 77.260556109, 4.9117755899, 96.6638761017, 96.7105583936, 86.773391397, 49.5325371648};
test_label[3371] = '{86.773391397};
test_output[3371] = '{10.6072701486};
############ END DEBUG ############*/
test_input[26976:26983] = '{32'hc2256fc6, 32'h42b28839, 32'hc0c42d6d, 32'h42a044d3, 32'hc2c3d893, 32'h427f3db9, 32'hc25bb130, 32'hc2ad4189};
test_label[3372] = '{32'hc2ad4189};
test_output[3372] = '{32'h432fe4e8};
/*############ DEBUG ############
test_input[26976:26983] = '{-41.3591549653, 89.2660619209, -6.13054529557, 80.13442243, -97.9229962702, 63.8102768973, -54.9230353616, -86.628000091};
test_label[3372] = '{-86.628000091};
test_output[3372] = '{175.894170194};
############ END DEBUG ############*/
test_input[26984:26991] = '{32'h3f988b50, 32'h41e52cc4, 32'hc261e695, 32'h42c2f9df, 32'hc2bf5f0b, 32'hc2af7375, 32'h41fea9a6, 32'hc079d968};
test_label[3373] = '{32'h3f988b50};
test_output[3373] = '{32'h42c097b2};
/*############ DEBUG ############
test_input[26984:26991] = '{1.19175142486, 28.6468588519, -56.4751777598, 97.4880330918, -95.6856301421, -87.7255036536, 31.8328362913, -3.90389445612};
test_label[3373] = '{1.19175142486};
test_output[3373] = '{96.2962816669};
############ END DEBUG ############*/
test_input[26992:26999] = '{32'hc186826b, 32'hc2946e50, 32'hc109f8da, 32'h41d319f4, 32'hc270c326, 32'hc2b35739, 32'h429345f9, 32'hc1c50b6e};
test_label[3374] = '{32'h429345f9};
test_output[3374] = '{32'h80000000};
/*############ DEBUG ############
test_input[26992:26999] = '{-16.8136799527, -74.2154548374, -8.62325473237, 26.3876722312, -60.1905730676, -89.6703592165, 73.6366648339, -24.630581527};
test_label[3374] = '{73.6366648339};
test_output[3374] = '{-0.0};
############ END DEBUG ############*/
test_input[27000:27007] = '{32'hc2900cd3, 32'h41f47176, 32'h42b1b754, 32'h428f91a8, 32'h42ac802b, 32'hc299bfed, 32'h428b0cdd, 32'h42189342};
test_label[3375] = '{32'h42b1b754};
test_output[3375] = '{32'h3d91a34d};
/*############ DEBUG ############
test_input[27000:27007] = '{-72.0250506669, 30.5554012951, 88.8580600435, 71.7844883269, 86.25033066, -76.8748539996, 69.5251250979, 38.1438064584};
test_label[3375] = '{88.8580600435};
test_output[3375] = '{0.0711122523902};
############ END DEBUG ############*/
test_input[27008:27015] = '{32'h428916c2, 32'h4282354d, 32'h4286d3a7, 32'hc2a292d9, 32'h42bd7b67, 32'hc29c3c96, 32'h42b7d9c8, 32'h42b6a64d};
test_label[3376] = '{32'hc29c3c96};
test_output[3376] = '{32'h432cf2b0};
/*############ DEBUG ############
test_input[27008:27015] = '{68.5444452006, 65.1041027707, 67.4133854301, -81.2868112112, 94.741018318, -78.1183326114, 91.9253552733, 91.3248030382};
test_label[3376] = '{-78.1183326114};
test_output[3376] = '{172.94800399};
############ END DEBUG ############*/
test_input[27016:27023] = '{32'hc2b5a25e, 32'h42ba6aed, 32'hc220c062, 32'h42020bab, 32'hc28a9405, 32'h41e38c4c, 32'h42c4a7a0, 32'hc164a2a7};
test_label[3377] = '{32'hc164a2a7};
test_output[3377] = '{32'h42e13f03};
/*############ DEBUG ############
test_input[27016:27023] = '{-90.8171228224, 93.2088359774, -40.1878744691, 32.511395412, -69.2891024694, 28.4435047137, 98.3273956898, -14.2897100969};
test_label[3377] = '{-14.2897100969};
test_output[3377] = '{112.623072586};
############ END DEBUG ############*/
test_input[27024:27031] = '{32'hc293d448, 32'hc28045e7, 32'hc194adde, 32'h40acc530, 32'h42227bc9, 32'h41137636, 32'hc252b487, 32'hc293bae9};
test_label[3378] = '{32'hc252b487};
test_output[3378] = '{32'h42ba9828};
/*############ DEBUG ############
test_input[27024:27031] = '{-73.9146108525, -64.1365262178, -18.5848954689, 5.39907079107, 40.6208833832, 9.21635990806, -52.6762945886, -73.8650586501};
test_label[3378] = '{-52.6762945886};
test_output[3378] = '{93.2971779719};
############ END DEBUG ############*/
test_input[27032:27039] = '{32'h428720a8, 32'h4184a988, 32'h42bd4ec7, 32'hc2a31755, 32'h413e294b, 32'hc21a4a3d, 32'h421d1844, 32'hc2296d1f};
test_label[3379] = '{32'hc21a4a3d};
test_output[3379] = '{32'h430539f3};
/*############ DEBUG ############
test_input[27032:27039] = '{67.5637805679, 16.5827782894, 94.6538596869, -81.5455675025, 11.8850814161, -38.5725002252, 39.2736958051, -42.3565651349};
test_label[3379] = '{-38.5725002252};
test_output[3379] = '{133.226359912};
############ END DEBUG ############*/
test_input[27040:27047] = '{32'h4276482e, 32'hc287d2b9, 32'hc2334a57, 32'h4271f357, 32'hc2a828ca, 32'hc18170f7, 32'hc251e529, 32'h42808082};
test_label[3380] = '{32'h4276482e};
test_output[3380] = '{32'h40312b61};
/*############ DEBUG ############
test_input[27040:27047] = '{61.5704868393, -67.9115708236, -44.822597286, 60.4876373333, -84.079668208, -16.1801582317, -52.4737875811, 64.2509919976};
test_label[3380] = '{61.5704868393};
test_output[3380] = '{2.76827268168};
############ END DEBUG ############*/
test_input[27048:27055] = '{32'h42b8da7e, 32'h41f6a95a, 32'hc2510ece, 32'h42b6a965, 32'hc24bf1b1, 32'h4261e827, 32'h419e5f3c, 32'hc1af2a68};
test_label[3381] = '{32'h419e5f3c};
test_output[3381] = '{32'h4291d653};
/*############ DEBUG ############
test_input[27048:27055] = '{92.4267392299, 30.8326915712, -52.2644581225, 91.33084997, -50.9860252121, 56.4767097413, 19.7965017311, -21.8957057783};
test_label[3381] = '{19.7965017311};
test_output[3381] = '{72.9186010239};
############ END DEBUG ############*/
test_input[27056:27063] = '{32'hc2b125b0, 32'hc1a7e830, 32'h42aa9c1c, 32'hc28eadb0, 32'hc2230899, 32'h41ff86c6, 32'hc0e4f2ab, 32'hc264859e};
test_label[3382] = '{32'hc264859e};
test_output[3382] = '{32'h430e6f75};
/*############ DEBUG ############
test_input[27056:27063] = '{-88.5736098076, -20.9883728224, 85.304900829, -71.3392337723, -40.7583944162, 31.940807822, -7.15462260457, -57.13048484};
test_label[3382] = '{-57.13048484};
test_output[3382] = '{142.435385669};
############ END DEBUG ############*/
test_input[27064:27071] = '{32'h4134e872, 32'hc203969c, 32'hc28c3c7b, 32'hc23658bd, 32'h42942da8, 32'h42014805, 32'hc21b6e90, 32'hc2c4943a};
test_label[3383] = '{32'h4134e872};
test_output[3383] = '{32'h427b2133};
/*############ DEBUG ############
test_input[27064:27071] = '{11.3067494483, -32.8970801052, -70.1181285355, -45.5866602919, 74.0891687844, 32.3203299287, -38.8579711748, -98.2895083393};
test_label[3383] = '{11.3067494483};
test_output[3383] = '{62.7824193361};
############ END DEBUG ############*/
test_input[27072:27079] = '{32'h42c3fc29, 32'hc24e928e, 32'hc2b406f3, 32'h41b4e6e2, 32'hc241e199, 32'h42b06438, 32'h40970d2e, 32'hc2be4744};
test_label[3384] = '{32'hc241e199};
test_output[3384] = '{32'h4312767f};
/*############ DEBUG ############
test_input[27072:27079] = '{97.9925034922, -51.6431214787, -90.0135726984, 22.6127349204, -48.4703117678, 88.1957421844, 4.72035899564, -95.1391936419};
test_label[3384] = '{-48.4703117678};
test_output[3384] = '{146.46287089};
############ END DEBUG ############*/
test_input[27080:27087] = '{32'h42b7a7b5, 32'h42afae39, 32'hbf4edfb6, 32'hc29b3ae7, 32'h42b98d8d, 32'h41d77515, 32'hc2850cb1, 32'hc28a21b9};
test_label[3385] = '{32'hc2850cb1};
test_output[3385] = '{32'h431fa239};
/*############ DEBUG ############
test_input[27080:27087] = '{91.8275515134, 87.8402758785, -0.808101048637, -77.6150423189, 92.7764685023, 26.9321686646, -66.5247903705, -69.0658647605};
test_label[3385] = '{-66.5247903705};
test_output[3385] = '{159.633681482};
############ END DEBUG ############*/
test_input[27088:27095] = '{32'hc22aaf1e, 32'hc03b9fcd, 32'h41f82859, 32'h42bc2318, 32'hc0d864e6, 32'h419891e3, 32'h429d9257, 32'hc2a08328};
test_label[3386] = '{32'h429d9257};
test_output[3386] = '{32'h41748609};
/*############ DEBUG ############
test_input[27088:27095] = '{-42.6710141029, -2.9316285342, 31.0197005366, 94.0685431258, -6.76231649888, 19.0712333562, 78.7858199122, -80.2561676619};
test_label[3386] = '{78.7858199122};
test_output[3386] = '{15.2827234442};
############ END DEBUG ############*/
test_input[27096:27103] = '{32'h42c14c9f, 32'hc1d40bf1, 32'hc1464814, 32'h4195bc2c, 32'hc27db017, 32'h420885b6, 32'hc2982182, 32'hc0dc2357};
test_label[3387] = '{32'hc27db017};
test_output[3387] = '{32'h43201255};
/*############ DEBUG ############
test_input[27096:27103] = '{96.649648268, -26.505831135, -12.3925973387, 18.716881153, -63.4219620054, 34.1305777205, -76.0654487276, -6.87931376206};
test_label[3387] = '{-63.4219620054};
test_output[3387] = '{160.071610273};
############ END DEBUG ############*/
test_input[27104:27111] = '{32'h42864ccb, 32'h41c7e341, 32'hc2833d1e, 32'h42c432ff, 32'h424589b1, 32'hc1ca9ce2, 32'h4296a038, 32'hc1a237e9};
test_label[3388] = '{32'h41c7e341};
test_output[3388] = '{32'h42923a2f};
/*############ DEBUG ############
test_input[27104:27111] = '{67.1499896322, 24.9859630707, -65.6193657829, 98.0996046039, 49.3844647458, -25.326602768, 75.3129273269, -20.2773007668};
test_label[3388] = '{24.9859630707};
test_output[3388] = '{73.1136415333};
############ END DEBUG ############*/
test_input[27112:27119] = '{32'hc25f9bd7, 32'h42532ff6, 32'hc1437cfd, 32'hc283e076, 32'h41260436, 32'h4272281b, 32'hc261fbd2, 32'hc224538d};
test_label[3389] = '{32'hc224538d};
test_output[3389] = '{32'h42cb3e0d};
/*############ DEBUG ############
test_input[27112:27119] = '{-55.9021889563, 52.7968382776, -12.2180149542, -65.9384040101, 10.3760283981, 60.5391652649, -56.4959190609, -41.0815910448};
test_label[3389] = '{-41.0815910448};
test_output[3389] = '{101.621190276};
############ END DEBUG ############*/
test_input[27120:27127] = '{32'hc1f5b8a3, 32'h42155c2a, 32'h429f46dc, 32'h42167188, 32'h424cc01c, 32'h4245d940, 32'hc1613886, 32'h4239a38c};
test_label[3390] = '{32'h429f46dc};
test_output[3390] = '{32'h2b132000};
/*############ DEBUG ############
test_input[27120:27127] = '{-30.715154451, 37.3400037483, 79.6383984524, 37.6108685925, 51.1876085223, 49.4621591355, -14.0762999454, 46.4097139578};
test_label[3390] = '{79.6383984524};
test_output[3390] = '{5.22692999994e-13};
############ END DEBUG ############*/
test_input[27128:27135] = '{32'h424653b9, 32'h42a73088, 32'hc12dbabe, 32'hc1ca482d, 32'h427592c8, 32'hc0af4143, 32'hc21cd0e8, 32'h4098f5ab};
test_label[3391] = '{32'hc12dbabe};
test_output[3391] = '{32'h42bce7df};
/*############ DEBUG ############
test_input[27128:27135] = '{49.5817595858, 83.594784316, -10.8580917146, -25.2852428876, 61.3933399182, -5.47671667929, -39.2040082941, 4.77998855217};
test_label[3391] = '{-10.8580917146};
test_output[3391] = '{94.4528760308};
############ END DEBUG ############*/
test_input[27136:27143] = '{32'h42baaf1a, 32'hc11fbfc7, 32'hc1da603b, 32'h42be8615, 32'h4277ab7e, 32'h4294d83f, 32'hc1e2a281, 32'hc1c3d7b1};
test_label[3392] = '{32'hc1da603b};
test_output[3392] = '{32'h42f56431};
/*############ DEBUG ############
test_input[27136:27143] = '{93.3419972026, -9.98432101718, -27.29698787, 95.2618790385, 61.9174741645, 74.4223535193, -28.3293477959, -24.4803175585};
test_label[3392] = '{-27.29698787};
test_output[3392] = '{122.695689132};
############ END DEBUG ############*/
test_input[27144:27151] = '{32'hc2595867, 32'h429cbd11, 32'h423b4bde, 32'hc29015b1, 32'hc0d93e4d, 32'hc22fe15a, 32'h42944956, 32'hc2346b09};
test_label[3393] = '{32'hc2595867};
test_output[3393] = '{32'h4304b859};
/*############ DEBUG ############
test_input[27144:27151] = '{-54.3363319363, 78.3692728511, 46.8240906032, -72.0423665397, -6.78885490163, -43.970071119, 74.1432376962, -45.1045281783};
test_label[3393] = '{-54.3363319363};
test_output[3393] = '{132.72010929};
############ END DEBUG ############*/
test_input[27152:27159] = '{32'h41c6c509, 32'h42c77eda, 32'hc1aa5e5e, 32'hc186199d, 32'h42a17213, 32'hc24eeea4, 32'h42882127, 32'h4284bb2d};
test_label[3394] = '{32'h42882127};
test_output[3394] = '{32'h41fd76cd};
/*############ DEBUG ############
test_input[27152:27159] = '{24.846209221, 99.7477588719, -21.2960774642, -16.7625055943, 80.7228036146, -51.7330457782, 68.0647511951, 66.3655778678};
test_label[3394] = '{68.0647511951};
test_output[3394] = '{31.6830076823};
############ END DEBUG ############*/
test_input[27160:27167] = '{32'hc2871d9b, 32'h4200c7b9, 32'h4209d2ae, 32'h41df5660, 32'h41097636, 32'hc2b66cf3, 32'hc213b389, 32'hc2a2e63e};
test_label[3395] = '{32'h41097636};
test_output[3395] = '{32'h41cfb814};
/*############ DEBUG ############
test_input[27160:27167] = '{-67.5578253636, 32.1950398054, 34.4557417911, 27.9171748879, 8.59136047494, -91.212789147, -36.9253288161, -81.449690536};
test_label[3395] = '{8.59136047494};
test_output[3395] = '{25.9648814756};
############ END DEBUG ############*/
test_input[27168:27175] = '{32'hc25c5446, 32'hc2c0645b, 32'hc2c72efc, 32'h41da1adb, 32'hc203e24e, 32'h42b56720, 32'hc2552f32, 32'h419378f2};
test_label[3396] = '{32'hc2c0645b};
test_output[3396] = '{32'h433ae5bd};
/*############ DEBUG ############
test_input[27168:27175] = '{-55.0822997609, -96.1960032235, -99.5917679647, 27.2631134892, -32.9710013627, 90.7014134214, -53.2960888876, 18.4340551093};
test_label[3396] = '{-96.1960032235};
test_output[3396] = '{186.897416645};
############ END DEBUG ############*/
test_input[27176:27183] = '{32'hc2b75548, 32'hc2b77341, 32'hbf1f8ff9, 32'h42a59604, 32'hc281d204, 32'hc2703843, 32'hc2a9f05a, 32'hc24ec7de};
test_label[3397] = '{32'hc24ec7de};
test_output[3397] = '{32'h43067cf9};
/*############ DEBUG ############
test_input[27176:27183] = '{-91.6665614712, -91.7251064557, -0.623290591886, 82.7929970329, -64.9101905322, -60.0549414996, -84.9694359827, -51.695182224};
test_label[3397] = '{-51.695182224};
test_output[3397] = '{134.488179257};
############ END DEBUG ############*/
test_input[27184:27191] = '{32'hc0fdc7e3, 32'h423beac9, 32'h4293e84a, 32'hc2a73246, 32'hc221acc9, 32'h40b06fe4, 32'hc094dfb3, 32'h413331fb};
test_label[3398] = '{32'h423beac9};
test_output[3398] = '{32'h41d7cb99};
/*############ DEBUG ############
test_input[27184:27191] = '{-7.9306501176, 46.9792808234, 73.9536929376, -83.5981908343, -40.4187342615, 5.51365861295, -4.6523070689, 11.1997019612};
test_label[3398] = '{46.9792808234};
test_output[3398] = '{26.9744121142};
############ END DEBUG ############*/
test_input[27192:27199] = '{32'h42b400f2, 32'hc25f9069, 32'h4201fa3e, 32'h4296609a, 32'h4292427b, 32'hc2649916, 32'hc2130659, 32'hc2a2f812};
test_label[3399] = '{32'h4296609a};
test_output[3399] = '{32'h416d02bc};
/*############ DEBUG ############
test_input[27192:27199] = '{90.0018442639, -55.8910246289, 32.4943788137, 75.1886771447, 73.1298415375, -57.1494961564, -36.7561984726, -81.48450961};
test_label[3399] = '{75.1886771447};
test_output[3399] = '{14.8131675351};
############ END DEBUG ############*/
test_input[27200:27207] = '{32'hc25bf800, 32'h4240e62a, 32'hc27d618d, 32'hc0f37eb5, 32'hc1d68ec6, 32'h423274de, 32'hc1c7116c, 32'h42a1255d};
test_label[3400] = '{32'hc1c7116c};
test_output[3400] = '{32'h42d2e9b8};
/*############ DEBUG ############
test_input[27200:27207] = '{-54.9921864129, 48.2247709065, -63.3452634553, -7.60921732035, -26.8197142108, 44.6141284187, -24.8835076991, 80.5729715414};
test_label[3400] = '{-24.8835076991};
test_output[3400] = '{105.45647924};
############ END DEBUG ############*/
test_input[27208:27215] = '{32'h41069c18, 32'h4261c776, 32'h40f51705, 32'hc269bcef, 32'h42bbdbaa, 32'h41eccfcc, 32'h4215d396, 32'hc23c6584};
test_label[3401] = '{32'h42bbdbaa};
test_output[3401] = '{32'h80000000};
/*############ DEBUG ############
test_input[27208:27215] = '{8.41310925869, 56.4447843308, 7.65906014622, -58.4345073624, 93.9290279831, 29.6014639985, 37.4566255151, -47.0991359651};
test_label[3401] = '{93.9290279831};
test_output[3401] = '{-0.0};
############ END DEBUG ############*/
test_input[27216:27223] = '{32'h42ad9a65, 32'hc1bfd0b2, 32'h42c5401e, 32'hc02fd5b5, 32'hc12d1763, 32'h42b70e6c, 32'h428e8181, 32'hc2c642a7};
test_label[3402] = '{32'hc02fd5b5};
test_output[3402] = '{32'h42cabf39};
/*############ DEBUG ############
test_input[27216:27223] = '{86.8015553719, -23.9769012125, 98.6252289709, -2.74741867321, -10.818209659, 91.5281658831, 71.2529351621, -99.1301836755};
test_label[3402] = '{-2.74741867321};
test_output[3402] = '{101.373482157};
############ END DEBUG ############*/
test_input[27224:27231] = '{32'h41ead4bf, 32'h419c10e4, 32'h41f2593e, 32'h4235b70a, 32'h40f4967d, 32'h422010b1, 32'h42863668, 32'h4238bbcf};
test_label[3403] = '{32'h419c10e4};
test_output[3403] = '{32'h423e645d};
/*############ DEBUG ############
test_input[27224:27231] = '{29.3538805951, 19.5082464492, 30.2935758025, 45.428747514, 7.6433703754, 40.0162990938, 67.1062588969, 46.1834049478};
test_label[3403] = '{19.5082464492};
test_output[3403] = '{47.5980124489};
############ END DEBUG ############*/
test_input[27232:27239] = '{32'h42a7e151, 32'h42bdec53, 32'h3f4e1c11, 32'h41e86481, 32'hc28a4ceb, 32'h40630066, 32'hc295d384, 32'h423183f5};
test_label[3404] = '{32'hc295d384};
test_output[3404] = '{32'h4329dfec};
/*############ DEBUG ############
test_input[27232:27239] = '{83.9400733296, 94.9615699707, 0.805115778201, 29.0490737499, -69.1502307855, 3.54689935437, -74.9131138995, 44.3788625775};
test_label[3404] = '{-74.9131138995};
test_output[3404] = '{169.874700217};
############ END DEBUG ############*/
test_input[27240:27247] = '{32'hc2b8496b, 32'h4266b7f9, 32'h42c4570d, 32'hc2277c46, 32'hc2086764, 32'hc22e9a08, 32'h410892d0, 32'hc25ee808};
test_label[3405] = '{32'h4266b7f9};
test_output[3405] = '{32'h4221f621};
/*############ DEBUG ############
test_input[27240:27247] = '{-92.1433980468, 57.6796591368, 98.1700205861, -41.8713611384, -34.100969187, -43.6504226387, 8.53584286411, -55.726593417};
test_label[3405] = '{57.6796591368};
test_output[3405] = '{40.4903614493};
############ END DEBUG ############*/
test_input[27248:27255] = '{32'h426f3121, 32'hc26cfbf3, 32'hc27a1b6c, 32'hc2418339, 32'hc1f33a53, 32'hc20c0de6, 32'h422b40b5, 32'h429c4f6f};
test_label[3406] = '{32'h426f3121};
test_output[3406] = '{32'h4192db7c};
/*############ DEBUG ############
test_input[27248:27255] = '{59.797976331, -59.2460452048, -62.5267789269, -48.3781487578, -30.4034788156, -35.01357364, 42.8131886127, 78.155145878};
test_label[3406] = '{59.797976331};
test_output[3406] = '{18.3571695577};
############ END DEBUG ############*/
test_input[27256:27263] = '{32'hc18ff05d, 32'h42bacb85, 32'h424391b9, 32'hc2a2de30, 32'h4209600b, 32'hc25eb9cf, 32'h41f4098e, 32'hc298a82b};
test_label[3407] = '{32'h42bacb85};
test_output[3407] = '{32'h80000000};
/*############ DEBUG ############
test_input[27256:27263] = '{-17.9923640747, 93.3975012781, 48.8923062124, -81.4339575846, 34.3437925834, -55.6814535126, 30.5046649707, -76.3284540383};
test_label[3407] = '{93.3975012781};
test_output[3407] = '{-0.0};
############ END DEBUG ############*/
test_input[27264:27271] = '{32'hc14ff747, 32'hc2c3a60d, 32'hc2ad4e96, 32'h404e8486, 32'h410191bf, 32'h41ca2584, 32'h4237e436, 32'hc24f08ff};
test_label[3408] = '{32'hc2c3a60d};
test_output[3408] = '{32'h430fcc14};
/*############ DEBUG ############
test_input[27264:27271] = '{-12.9978706227, -97.8243209684, -86.6534916773, 3.22683860253, 8.09808230516, 25.2683191129, 45.9728627042, -51.7587837657};
test_label[3408] = '{-97.8243209684};
test_output[3408] = '{143.797183674};
############ END DEBUG ############*/
test_input[27272:27279] = '{32'hc1b6d3f2, 32'hc2022653, 32'hc13d5fbb, 32'h4246dba6, 32'h42986058, 32'h42c14cdd, 32'h42b7b0be, 32'hc1e768dc};
test_label[3409] = '{32'hc13d5fbb};
test_output[3409] = '{32'h42d8fd01};
/*############ DEBUG ############
test_input[27272:27279] = '{-22.8534888144, -32.5374249162, -11.835871242, 49.7145017456, 76.1881691727, 96.6501239004, 91.8451999641, -28.9262012435};
test_label[3409] = '{-11.835871242};
test_output[3409] = '{108.494151117};
############ END DEBUG ############*/
test_input[27280:27287] = '{32'h41fe0cef, 32'h428c8ebc, 32'hc186b0de, 32'h412dcb81, 32'h421f3831, 32'hc2b86287, 32'h4250ce7a, 32'h425f512e};
test_label[3410] = '{32'hc2b86287};
test_output[3410] = '{32'h432278a2};
/*############ DEBUG ############
test_input[27280:27287] = '{31.756315024, 70.2787747468, -16.8363612883, 10.8621838262, 39.8048759454, -92.1924399562, 52.2016373468, 55.8292772415};
test_label[3410] = '{-92.1924399562};
test_output[3410] = '{162.471215248};
############ END DEBUG ############*/
test_input[27288:27295] = '{32'hc2be20e2, 32'hc17672f7, 32'h41fd9808, 32'h42bd9674, 32'h40c1deab, 32'h42a24381, 32'h415e8b83, 32'h42118c70};
test_label[3411] = '{32'h41fd9808};
test_output[3411] = '{32'h427c60e4};
/*############ DEBUG ############
test_input[27288:27295] = '{-95.0642251412, -15.4030671331, 31.6992334537, 94.7938520986, 6.05843102585, 81.1318447696, 13.909060259, 36.3871446784};
test_label[3411] = '{31.6992334537};
test_output[3411] = '{63.0946198108};
############ END DEBUG ############*/
test_input[27296:27303] = '{32'hc2bc61a1, 32'h4224d0be, 32'h42a9d18a, 32'hc1ccd552, 32'hc212783f, 32'h417da573, 32'hc1b32e7b, 32'h428db621};
test_label[3412] = '{32'hc1ccd552};
test_output[3412] = '{32'h42dd06df};
/*############ DEBUG ############
test_input[27296:27303] = '{-94.1906832777, 41.2038481438, 84.9092584981, -25.6041600747, -36.6174293388, 15.852892832, -22.3976963499, 70.8557214088};
test_label[3412] = '{-25.6041600747};
test_output[3412] = '{110.513419361};
############ END DEBUG ############*/
test_input[27304:27311] = '{32'h429e8af9, 32'hc13dbfbb, 32'hc2217ef4, 32'hc20a9bba, 32'hc1b8fbd4, 32'hc24e47a5, 32'hc1e25a91, 32'hc25b474b};
test_label[3413] = '{32'hc1e25a91};
test_output[3413] = '{32'h42d7219d};
/*############ DEBUG ############
test_input[27304:27311] = '{79.2714306903, -11.8593093171, -40.3739778718, -34.6520753, -23.1229628742, -51.569964069, -28.294221475, -54.8196208723};
test_label[3413] = '{-28.294221475};
test_output[3413] = '{107.565652165};
############ END DEBUG ############*/
test_input[27312:27319] = '{32'h427958d5, 32'hc290e51a, 32'h41c1ed81, 32'hc29a66c8, 32'hc181999e, 32'hc1b41a67, 32'hc219b426, 32'h42a03ba0};
test_label[3414] = '{32'hc219b426};
test_output[3414] = '{32'h42ed15b3};
/*############ DEBUG ############
test_input[27312:27319] = '{62.336750647, -72.4474675855, 24.2409688095, -77.2007417667, -16.2000077212, -22.5128913016, -38.4259258393, 80.1164543764};
test_label[3414] = '{-38.4259258393};
test_output[3414] = '{118.542380235};
############ END DEBUG ############*/
test_input[27320:27327] = '{32'h4261daaf, 32'h41e39e35, 32'h42883dd7, 32'hc1956288, 32'h4102296f, 32'h42a450d5, 32'h4293e749, 32'h42c1bb5b};
test_label[3415] = '{32'h4261daaf};
test_output[3415] = '{32'h42219c06};
/*############ DEBUG ############
test_input[27320:27327] = '{56.4635586449, 28.4522493888, 68.1207826426, -18.6731108274, 8.135115236, 82.1578752013, 73.9517271836, 96.8659251235};
test_label[3415] = '{56.4635586449};
test_output[3415] = '{40.4023668883};
############ END DEBUG ############*/
test_input[27328:27335] = '{32'hc19a379f, 32'hc1267b07, 32'h426f7f4b, 32'hc1345e5f, 32'hc2932230, 32'hc28e853b, 32'hc21d8fcd, 32'hc287f741};
test_label[3416] = '{32'hc19a379f};
test_output[3416] = '{32'h429e4d8d};
/*############ DEBUG ############
test_input[27328:27335] = '{-19.2771583975, -10.4050355302, 59.8743103079, -11.273040118, -73.5667692006, -71.2602129194, -39.3904304228, -67.9829192686};
test_label[3416] = '{-19.2771583975};
test_output[3416] = '{79.1514687054};
############ END DEBUG ############*/
test_input[27336:27343] = '{32'hc26f370e, 32'hc2ab4e14, 32'hc2ad4cee, 32'h42a775fa, 32'hc1ab0814, 32'h42a1ef96, 32'h428aeff0, 32'hc09ae8ba};
test_label[3417] = '{32'h42a1ef96};
test_output[3417] = '{32'h4034b789};
/*############ DEBUG ############
test_input[27336:27343] = '{-59.8037647375, -85.6524959185, -86.6502523896, 83.7304202246, -21.3789439221, 80.967940917, 69.4686307632, -4.84090920729};
test_label[3417] = '{80.967940917};
test_output[3417] = '{2.82370204041};
############ END DEBUG ############*/
test_input[27344:27351] = '{32'hc27c5b02, 32'h42231639, 32'h429e9401, 32'hc1584fbf, 32'hc29a4682, 32'h424807c0, 32'hc1a35044, 32'h427a8739};
test_label[3418] = '{32'h429e9401};
test_output[3418] = '{32'h337a8f19};
/*############ DEBUG ############
test_input[27344:27351] = '{-63.0888756794, 40.771702536, 79.2890722712, -13.5194692243, -77.1377140073, 50.0075702027, -20.4141920426, 62.6320535635};
test_label[3418] = '{79.2890722712};
test_output[3418] = '{5.83378079541e-08};
############ END DEBUG ############*/
test_input[27352:27359] = '{32'h41a49899, 32'h42a811f7, 32'hc22bef5b, 32'h422732da, 32'hc1b05943, 32'hc2120d98, 32'hc022e70b, 32'hc2a113c0};
test_label[3419] = '{32'hc2a113c0};
test_output[3419] = '{32'h432492dc};
/*############ DEBUG ############
test_input[27352:27359] = '{20.5745097737, 84.0350904122, -42.9837472419, 41.799660899, -22.0435839486, -36.5132736486, -2.5453516439, -80.5385761642};
test_label[3419] = '{-80.5385761642};
test_output[3419] = '{164.573666576};
############ END DEBUG ############*/
test_input[27360:27367] = '{32'h4231d0da, 32'h425366d1, 32'h3fb75c79, 32'h42b00b92, 32'h421f5b08, 32'hc2803dab, 32'h421f7f3a, 32'hc2aef758};
test_label[3420] = '{32'h421f5b08};
test_output[3420] = '{32'h4240bc1c};
/*############ DEBUG ############
test_input[27360:27367] = '{44.4539560652, 52.8504056225, 1.43250951526, 88.0225996712, 39.8388974831, -64.1204417939, 39.8742431551, -87.4830965965};
test_label[3420] = '{39.8388974831};
test_output[3420] = '{48.1837021881};
############ END DEBUG ############*/
test_input[27368:27375] = '{32'h41b34fff, 32'hc1adda1b, 32'h411d43a9, 32'h42b8cf27, 32'hc1daf427, 32'h42a7320b, 32'h41f4e702, 32'h428a8cc9};
test_label[3421] = '{32'h41f4e702};
test_output[3421] = '{32'h42772af5};
/*############ DEBUG ############
test_input[27368:27375] = '{22.414059804, -21.7314960913, 9.82901827145, 92.4045971017, -27.3692159543, 83.5977381939, 30.6127966506, 69.274969517};
test_label[3421] = '{30.6127966506};
test_output[3421] = '{61.7919501428};
############ END DEBUG ############*/
test_input[27376:27383] = '{32'h410db498, 32'h42a3ca13, 32'h41bd69e7, 32'h42c76fdd, 32'hc1046065, 32'h405adf74, 32'h4207feb2, 32'hc216bef7};
test_label[3422] = '{32'h42c76fdd};
test_output[3422] = '{32'h329c07a1};
/*############ DEBUG ############
test_input[27376:27383] = '{8.85659043787, 81.894676638, 23.6767094046, 99.7184865781, -8.27353387686, 3.41988839433, 33.9987243636, -37.6864885062};
test_label[3422] = '{99.7184865781};
test_output[3422] = '{1.81642593728e-08};
############ END DEBUG ############*/
test_input[27384:27391] = '{32'hc29ded89, 32'hc2364a5f, 32'h421493d1, 32'h420cf5aa, 32'hc2889a61, 32'hc2a36441, 32'hc2c4ebd9, 32'h42bc3cca};
test_label[3423] = '{32'hc29ded89};
test_output[3423] = '{32'h432d152a};
/*############ DEBUG ############
test_input[27384:27391] = '{-78.9639388302, -45.5726277089, 37.1443513377, 35.2399048741, -68.3015216798, -81.6958057555, -98.4606362954, 94.1187309576};
test_label[3423] = '{-78.9639388302};
test_output[3423] = '{173.082669788};
############ END DEBUG ############*/
test_input[27392:27399] = '{32'h42c314d8, 32'h4260c268, 32'hc20a65c8, 32'hc1a1b1c9, 32'h416b07aa, 32'hc1da5aa6, 32'h42588000, 32'h41732a17};
test_label[3424] = '{32'h416b07aa};
test_output[3424] = '{32'h42a5b3e2};
/*############ DEBUG ############
test_input[27392:27399] = '{97.5407071213, 56.1898494831, -34.5993955803, -20.2118083853, 14.6893708235, -27.2942618209, 54.1249998705, 15.1977755857};
test_label[3424] = '{14.6893708235};
test_output[3424] = '{82.8513362978};
############ END DEBUG ############*/
test_input[27400:27407] = '{32'hc2c04850, 32'hc2b647fc, 32'hc2639df7, 32'hc1653375, 32'h419995bf, 32'h41df3c43, 32'hc2272dff, 32'hc281a7a5};
test_label[3425] = '{32'hc1653375};
test_output[3425] = '{32'h4228eb2a};
/*############ DEBUG ############
test_input[27400:27407] = '{-96.1412353571, -91.1405920264, -56.9042635176, -14.3250625178, 19.1981174724, 27.9044252553, -41.7949168381, -64.8274298841};
test_label[3425] = '{-14.3250625178};
test_output[3425] = '{42.2296532977};
############ END DEBUG ############*/
test_input[27408:27415] = '{32'hc205bec6, 32'h41fde8f4, 32'hc2aca5a7, 32'hc237bbf6, 32'h42699d81, 32'hc2128b1b, 32'h42249809, 32'hc2a73483};
test_label[3426] = '{32'hc2128b1b};
test_output[3426] = '{32'h42be144e};
/*############ DEBUG ############
test_input[27408:27415] = '{-33.4363012447, 31.7387459564, -86.3235374035, -45.933555154, 58.4038111869, -36.6358464744, 41.1484717459, -83.6025587672};
test_label[3426] = '{-36.6358464744};
test_output[3426] = '{95.0396576934};
############ END DEBUG ############*/
test_input[27416:27423] = '{32'hc2485ed5, 32'hc22c6b5e, 32'h41507957, 32'hc16ab094, 32'hc1c7a548, 32'hc1b1e421, 32'h4244193d, 32'h42a12b1f};
test_label[3427] = '{32'hc1c7a548};
test_output[3427] = '{32'h42d31471};
/*############ DEBUG ############
test_input[27416:27423] = '{-50.0926080903, -43.1048490807, 13.0296240579, -14.6681094997, -24.9557028516, -22.236390816, 49.0246484473, 80.5842189963};
test_label[3427] = '{-24.9557028516};
test_output[3427] = '{105.539921848};
############ END DEBUG ############*/
test_input[27424:27431] = '{32'h42b306ad, 32'h42133788, 32'hc18524a1, 32'h41337cc5, 32'h41dd53fa, 32'hc1a76556, 32'h4231b1ac, 32'h42656c42};
test_label[3428] = '{32'hc18524a1};
test_output[3428] = '{32'h42d44fd5};
/*############ DEBUG ############
test_input[27424:27431] = '{89.5130407293, 36.8042300019, -16.6428843911, 11.2179611102, 27.6660042775, -20.9244796189, 44.4235064712, 57.3557219102};
test_label[3428] = '{-16.6428843911};
test_output[3428] = '{106.15592512};
############ END DEBUG ############*/
test_input[27432:27439] = '{32'h42c2d1d0, 32'h42bc41de, 32'h4023df1a, 32'hc2a73024, 32'hc155d5bb, 32'hc281ce8b, 32'hc2a69f90, 32'h424f2e0d};
test_label[3429] = '{32'hc281ce8b};
test_output[3429] = '{32'h432259a0};
/*############ DEBUG ############
test_input[27432:27439] = '{97.4097917071, 94.1286496773, 2.56049192057, -83.5940276505, -13.3646803469, -64.9034047081, -83.311645283, 51.7949722007};
test_label[3429] = '{-64.9034047081};
test_output[3429] = '{162.35009261};
############ END DEBUG ############*/
test_input[27440:27447] = '{32'h42c00722, 32'hc29539f2, 32'hc21ebe20, 32'hc2aa9f81, 32'hc28df298, 32'hc28601c2, 32'h41b34352, 32'h41a7ef23};
test_label[3430] = '{32'h41a7ef23};
test_output[3430] = '{32'h42960b59};
/*############ DEBUG ############
test_input[27440:27447] = '{96.0139319589, -74.6131758031, -39.6856688587, -85.311529661, -70.973816058, -67.0034300201, 22.4078703797, 20.9917659991};
test_label[3430] = '{20.9917659991};
test_output[3430] = '{75.0221659598};
############ END DEBUG ############*/
test_input[27448:27455] = '{32'h42b63a0d, 32'hc292f7a6, 32'hc251ff84, 32'h4109c633, 32'h41ff851c, 32'hc0e15828, 32'hc2c0e081, 32'hc0f1a9a3};
test_label[3431] = '{32'hc251ff84};
test_output[3431] = '{32'h430f9ce7};
/*############ DEBUG ############
test_input[27448:27455] = '{91.1133798479, -73.4836903575, -52.4995268055, 8.61088847667, 31.9399943151, -7.04201110072, -96.4384870736, -7.55195756619};
test_label[3431] = '{-52.4995268055};
test_output[3431] = '{143.612906653};
############ END DEBUG ############*/
test_input[27456:27463] = '{32'h4187e5e5, 32'hc27fa7ac, 32'hc2794b95, 32'h4003dfb5, 32'h422a0641, 32'hc2936efe, 32'hc28c346f, 32'h426cdc26};
test_label[3432] = '{32'h4003dfb5};
test_output[3432] = '{32'h42649e2b};
/*############ DEBUG ############
test_input[27456:27463] = '{16.9872536077, -63.9137424794, -62.3238088425, 2.06052902042, 42.506105999, -73.7167783661, -70.1024071113, 59.2149895365};
test_label[3432] = '{2.06052902042};
test_output[3432] = '{57.1544605715};
############ END DEBUG ############*/
test_input[27464:27471] = '{32'h4144ac75, 32'hc2c284ae, 32'h41d51d7a, 32'hc2bafa43, 32'h42b7154d, 32'hc2b691a1, 32'hc24ed438, 32'hc107c4d8};
test_label[3433] = '{32'hc2bafa43};
test_output[3433] = '{32'h433907c8};
/*############ DEBUG ############
test_input[27464:27471] = '{12.2921037462, -97.2591378307, 26.6393937133, -93.4887945288, 91.5416064408, -91.2844323955, -51.7072456797, -8.48555713572};
test_label[3433] = '{-93.4887945288};
test_output[3433] = '{185.03040097};
############ END DEBUG ############*/
test_input[27472:27479] = '{32'h421ce210, 32'hc1a946c7, 32'hc2878e2f, 32'h41dc971a, 32'h425dfad4, 32'hc2908841, 32'h428ecadd, 32'h42534519};
test_label[3434] = '{32'h425dfad4};
test_output[3434] = '{32'h417e6b95};
/*############ DEBUG ############
test_input[27472:27479] = '{39.2207649459, -21.1595593532, -67.7776998425, 27.5737797704, 55.4949491902, -72.2661226471, 71.3962138888, 52.8174767252};
test_label[3434] = '{55.4949491902};
test_output[3434] = '{15.9012648313};
############ END DEBUG ############*/
test_input[27480:27487] = '{32'h42bc8e22, 32'h429dfb6c, 32'hc228b28d, 32'h41f1614b, 32'h4086c92f, 32'h41d6c84e, 32'h40dc1d8c, 32'hc2a4efdb};
test_label[3435] = '{32'h41d6c84e};
test_output[3435] = '{32'h4286dc0f};
/*############ DEBUG ############
test_input[27480:27487] = '{94.2776049816, 78.9910571285, -42.1743655255, 30.1725064322, 4.21205875371, 26.8478043982, 6.87860684979, -82.4684711354};
test_label[3435] = '{26.8478043982};
test_output[3435] = '{67.4298008131};
############ END DEBUG ############*/
test_input[27488:27495] = '{32'h4251b4b0, 32'hc23037cf, 32'hc1efacf1, 32'hc22f958e, 32'h426026a7, 32'h41a7ac48, 32'hc138d041, 32'hc2b5bd3f};
test_label[3436] = '{32'hc138d041};
test_output[3436] = '{32'h42873b02};
/*############ DEBUG ############
test_input[27488:27495] = '{52.4264541673, -44.0545024445, -29.9594438095, -43.8960495464, 56.0377477861, 20.9591225169, -11.5508435017, -90.8696219623};
test_label[3436] = '{-11.5508435017};
test_output[3436] = '{67.6152496496};
############ END DEBUG ############*/
test_input[27496:27503] = '{32'hc1f40721, 32'hc1e26c47, 32'hc2b5648b, 32'h42c494b2, 32'hc2962d37, 32'hc23412ce, 32'h4208eb0f, 32'h4111849f};
test_label[3437] = '{32'hc1f40721};
test_output[3437] = '{32'h4300cb3d};
/*############ DEBUG ############
test_input[27496:27503] = '{-30.5034813823, -28.3028690093, -90.6963697151, 98.2904174198, -75.0883124125, -45.0183653692, 34.2295481895, 9.09487852212};
test_label[3437] = '{-30.5034813823};
test_output[3437] = '{128.793898802};
############ END DEBUG ############*/
test_input[27504:27511] = '{32'h42b606e6, 32'h4276fa48, 32'hc28d18a9, 32'h426b29ca, 32'h42b88f4c, 32'hc29a7aa3, 32'hc18ca885, 32'hc18f6668};
test_label[3438] = '{32'hc28d18a9};
test_output[3438] = '{32'h4323138b};
/*############ DEBUG ############
test_input[27504:27511] = '{91.013474267, 61.7444151613, -70.548167611, 58.7908097275, 92.2798781048, -77.2395273952, -17.5822844191, -17.9250024979};
test_label[3438] = '{-70.548167611};
test_output[3438] = '{163.07634488};
############ END DEBUG ############*/
test_input[27512:27519] = '{32'hc265a86b, 32'h4287d61c, 32'hc1a7b231, 32'h4229c740, 32'h421b3cf5, 32'h3fac6e47, 32'h424462d6, 32'hc2c04364};
test_label[3439] = '{32'hc265a86b};
test_output[3439] = '{32'h42faaa52};
/*############ DEBUG ############
test_input[27512:27519] = '{-57.4144713689, 67.9181832458, -20.9620077022, 42.4445792217, 38.8095282403, 1.34711537751, 49.0965207065, -96.1316204392};
test_label[3439] = '{-57.4144713689};
test_output[3439] = '{125.332654621};
############ END DEBUG ############*/
test_input[27520:27527] = '{32'hc201cb4b, 32'h4280d2b1, 32'h422c0266, 32'h4291de45, 32'h42bf9420, 32'h41b01ceb, 32'h42522afd, 32'h42a9abf8};
test_label[3440] = '{32'h42bf9420};
test_output[3440] = '{32'h3792c86c};
/*############ DEBUG ############
test_input[27520:27527] = '{-32.4485294101, 64.4115077465, 43.0023424724, 72.9341167728, 95.7893072642, 22.0141206992, 52.5419811213, 84.8358787281};
test_label[3440] = '{95.7893072642};
test_output[3440] = '{1.74978856323e-05};
############ END DEBUG ############*/
test_input[27528:27535] = '{32'hc2bf6581, 32'hc26c5641, 32'h41e7bb69, 32'hc214b3e2, 32'h42bad8f4, 32'h42b78c24, 32'h423a944f, 32'hc1db6dbf};
test_label[3441] = '{32'h42b78c24};
test_output[3441] = '{32'h3fe9b076};
/*############ DEBUG ############
test_input[27528:27535] = '{-95.6982515813, -59.0842340174, 28.966509316, -37.1756655093, 93.4237372373, 91.7737094974, 46.6448318112, -27.4285866222};
test_label[3441] = '{91.7737094974};
test_output[3441] = '{1.82569770822};
############ END DEBUG ############*/
test_input[27536:27543] = '{32'h42c1620b, 32'hc28049d9, 32'hc1ed72d1, 32'hc24c30dd, 32'hc13ee028, 32'h4167f144, 32'h4116a14c, 32'h4214df00};
test_label[3442] = '{32'h4214df00};
test_output[3442] = '{32'h426de516};
/*############ DEBUG ############
test_input[27536:27543] = '{96.6914902616, -64.1442345515, -29.6810633801, -51.0477193711, -11.9297254108, 14.4964027841, 9.4143792073, 37.2177725056};
test_label[3442] = '{37.2177725056};
test_output[3442] = '{59.473717756};
############ END DEBUG ############*/
test_input[27544:27551] = '{32'h41a0df9e, 32'h420fd520, 32'hc2504adf, 32'h41c9d409, 32'h408fb39d, 32'h41e266fe, 32'hc228917a, 32'hc1b35773};
test_label[3443] = '{32'hc228917a};
test_output[3443] = '{32'h429c338e};
/*############ DEBUG ############
test_input[27544:27551] = '{20.1091886561, 35.9581307242, -52.0731146254, 25.2285335401, 4.49067523053, 28.3002896098, -42.142067415, -22.4176994394};
test_label[3443] = '{-42.142067415};
test_output[3443] = '{78.1006923614};
############ END DEBUG ############*/
test_input[27552:27559] = '{32'h40221fa3, 32'hc239e758, 32'h41ac3d81, 32'h429102c9, 32'hc1ce0c50, 32'h4130a1e8, 32'h4202b47c, 32'hc18672e8};
test_label[3444] = '{32'hc18672e8};
test_output[3444] = '{32'h42b29f83};
/*############ DEBUG ############
test_input[27552:27559] = '{2.53318097161, -46.4759224613, 21.5300302568, 72.5054391306, -25.7560116144, 11.0395283094, 32.676252827, -16.8061065814};
test_label[3444] = '{-16.8061065814};
test_output[3444] = '{89.311545712};
############ END DEBUG ############*/
test_input[27560:27567] = '{32'h42586b51, 32'h41f3e98b, 32'h42c0361c, 32'h42be746b, 32'h42c7dd91, 32'h4200ce42, 32'hc2a98226, 32'hc285da3f};
test_label[3445] = '{32'h42c0361c};
test_output[3445] = '{32'h4076dfeb};
/*############ DEBUG ############
test_input[27560:27567] = '{54.1048005945, 30.4890350318, 96.1056846414, 95.2273798621, 99.9327467559, 32.2014240634, -84.7541936131, -66.9262646608};
test_label[3445] = '{96.1056846414};
test_output[3445] = '{3.8574167982};
############ END DEBUG ############*/
test_input[27568:27575] = '{32'hc159829c, 32'h410783b2, 32'hc2b656dc, 32'hc2c7a0ca, 32'h40b0ffe7, 32'hc2967de2, 32'h413a6af5, 32'h4269117f};
test_label[3446] = '{32'hc2967de2};
test_output[3446] = '{32'h43058351};
/*############ DEBUG ############
test_input[27568:27575] = '{-13.5943871627, 8.46965235349, -91.1696497296, -99.8140420302, 5.53123828117, -75.2458663536, 11.6511128479, 58.2670873836};
test_label[3446] = '{-75.2458663536};
test_output[3446] = '{133.512953737};
############ END DEBUG ############*/
test_input[27576:27583] = '{32'h422ab493, 32'h411dc114, 32'h42aff3a3, 32'h42a6d7d3, 32'hc2af8785, 32'h4286aced, 32'hc2a8157c, 32'h42957f90};
test_label[3447] = '{32'h42957f90};
test_output[3447] = '{32'h4153cb72};
/*############ DEBUG ############
test_input[27576:27583] = '{42.6763403163, 9.85963859546, 87.9758500568, 83.4215289022, -87.7646842324, 67.3377487363, -84.0419604474, 74.7491492092};
test_label[3447] = '{74.7491492092};
test_output[3447] = '{13.2371693049};
############ END DEBUG ############*/
test_input[27584:27591] = '{32'h41265610, 32'hc2bf8ad4, 32'h416f4d81, 32'hc039248e, 32'hc2c07aa1, 32'h423b3fb1, 32'h4201baf0, 32'hc2ad3a84};
test_label[3448] = '{32'h41265610};
test_output[3448] = '{32'h4211aa2d};
/*############ DEBUG ############
test_input[27584:27591] = '{10.3960114038, -95.7711477927, 14.9564222738, -2.89285609194, -96.2395115382, 46.8121987932, 32.4325574804, -86.6142921269};
test_label[3448] = '{10.3960114038};
test_output[3448] = '{36.4161879583};
############ END DEBUG ############*/
test_input[27592:27599] = '{32'h426c3575, 32'hc20b5b67, 32'hc24901e6, 32'h4282b6de, 32'hc28c3b9f, 32'h42b1dab8, 32'h41807f8b, 32'hc1d7818e};
test_label[3449] = '{32'h426c3575};
test_output[3449] = '{32'h41eefff8};
/*############ DEBUG ############
test_input[27592:27599] = '{59.0522022778, -34.8392592419, -50.251855129, 65.3571661541, -70.11644818, 88.9271860749, 16.0622777411, -26.938258339};
test_label[3449] = '{59.0522022778};
test_output[3449] = '{29.8749837972};
############ END DEBUG ############*/
test_input[27600:27607] = '{32'hc1f2839c, 32'hc23cd05c, 32'hc292d2d8, 32'hc180214d, 32'h426ba77d, 32'h42439c9f, 32'hc216fda1, 32'h420101f4};
test_label[3450] = '{32'hc23cd05c};
test_output[3450] = '{32'h42d43bf3};
/*############ DEBUG ############
test_input[27600:27607] = '{-30.3142621789, -47.2034754537, -73.4118035202, -16.016259782, 58.9135645162, 48.9029501596, -37.7476841678, 32.2519080744};
test_label[3450] = '{-47.2034754537};
test_output[3450] = '{106.11708489};
############ END DEBUG ############*/
test_input[27608:27615] = '{32'h428454c0, 32'h417334c6, 32'hc1b776e0, 32'hc2c4a47f, 32'h41745ffb, 32'h42965bc2, 32'h42474c0b, 32'h41f1e0b2};
test_label[3451] = '{32'h428454c0};
test_output[3451] = '{32'h41103892};
/*############ DEBUG ############
test_input[27608:27615] = '{66.1655260577, 15.2003843236, -22.9330446377, -98.3212795903, 15.2734326933, 75.1792157784, 49.8242603872, 30.2347153429};
test_label[3451] = '{66.1655260577};
test_output[3451] = '{9.01381144522};
############ END DEBUG ############*/
test_input[27616:27623] = '{32'h41d804d0, 32'h422c8dce, 32'hc29885e3, 32'h42b9eeec, 32'h423348d5, 32'h42c1f5fb, 32'hc261e015, 32'hc230a025};
test_label[3452] = '{32'h422c8dce};
test_output[3452] = '{32'h4257707e};
/*############ DEBUG ############
test_input[27616:27623] = '{27.0023505905, 43.1384815532, -76.2614966235, 92.9666460339, 44.8211242952, 96.9804319006, -56.4688295614, -44.1563927672};
test_label[3452] = '{43.1384815532};
test_output[3452] = '{53.8598539908};
############ END DEBUG ############*/
test_input[27624:27631] = '{32'h4020ebfe, 32'h42700214, 32'hc2a7b758, 32'h425ae866, 32'h427d3a64, 32'h4238ce2e, 32'hc2c6b1e1, 32'hc0ac1c7a};
test_label[3453] = '{32'hc2c6b1e1};
test_output[3453] = '{32'h4322b0cf};
/*############ DEBUG ############
test_input[27624:27631] = '{2.51440391269, 60.0020286988, -83.8580898253, 54.7269519729, 63.3070211395, 46.2013490702, -99.3474191916, -5.3784759092};
test_label[3453] = '{-99.3474191916};
test_output[3453] = '{162.690663613};
############ END DEBUG ############*/
test_input[27632:27639] = '{32'hc12845dc, 32'hc21af1db, 32'hc299cef6, 32'hc27735cd, 32'h424e5651, 32'h428671bd, 32'h422c586e, 32'h42937771};
test_label[3454] = '{32'h422c586e};
test_output[3454] = '{32'h41f52ff4};
/*############ DEBUG ############
test_input[27632:27639] = '{-10.5170550406, -38.7361886654, -76.9042239005, -61.8025413147, 51.584294803, 67.2221426793, 43.0863558545, 73.733285151};
test_label[3454] = '{43.0863558545};
test_output[3454] = '{30.6484149727};
############ END DEBUG ############*/
test_input[27640:27647] = '{32'h420b2df4, 32'hc24fdf37, 32'h411c9b8d, 32'hc18efb78, 32'h4146edc4, 32'hc2c29df5, 32'h427c0598, 32'h41b9ba04};
test_label[3455] = '{32'hc24fdf37};
test_output[3455] = '{32'h42e5f267};
/*############ DEBUG ############
test_input[27640:27647] = '{34.794875308, -51.9679839416, 9.78797656479, -17.8727876766, 12.4330481034, -97.3085086387, 63.0054608129, 23.2158284251};
test_label[3455] = '{-51.9679839416};
test_output[3455] = '{114.973444754};
############ END DEBUG ############*/
test_input[27648:27655] = '{32'h419565b2, 32'hc19938c5, 32'hc1cbc10c, 32'h427b92fe, 32'h41e2f5aa, 32'h42b44ec1, 32'h42ba8e20, 32'h41964c03};
test_label[3456] = '{32'hc19938c5};
test_output[3456] = '{32'h42e0f25c};
/*############ DEBUG ############
test_input[27648:27655] = '{18.6746552789, -19.1527185979, -25.4692608824, 62.8935482592, 28.369952798, 90.1538135359, 93.277584926, 18.7871156282};
test_label[3456] = '{-19.1527185979};
test_output[3456] = '{112.473354343};
############ END DEBUG ############*/
test_input[27656:27663] = '{32'h423bbe9b, 32'h429f1f2f, 32'hc2109de7, 32'h4189a0de, 32'h40d10e64, 32'h415a7184, 32'h4265a1eb, 32'hc24eaa92};
test_label[3457] = '{32'h4189a0de};
test_output[3457] = '{32'h42796def};
/*############ DEBUG ############
test_input[27656:27663] = '{46.936139821, 79.5609056435, -36.1542003336, 17.2035493308, 6.53300688137, 13.6527141642, 57.4081240647, -51.6665718667};
test_label[3457] = '{17.2035493308};
test_output[3457] = '{62.3573563129};
############ END DEBUG ############*/
test_input[27664:27671] = '{32'hc2341b82, 32'hc2bdc974, 32'h42ae9a9a, 32'h41a45f08, 32'h412ee720, 32'hc255c16b, 32'hc20ca974, 32'hc21f7289};
test_label[3458] = '{32'hc255c16b};
test_output[3458] = '{32'h430cbda8};
/*############ DEBUG ############
test_input[27664:27671] = '{-45.0268622236, -94.8934652725, 87.3019568599, 20.5464011159, 10.9314271416, -53.4388838965, -35.1654800116, -39.8618498155};
test_label[3458] = '{-53.4388838965};
test_output[3458] = '{140.740840756};
############ END DEBUG ############*/
test_input[27672:27679] = '{32'hc1ad6cb9, 32'h416d6d11, 32'hc259f12d, 32'hc1907764, 32'hc2a1691a, 32'h42468341, 32'h42957019, 32'hc2075001};
test_label[3459] = '{32'hc1ad6cb9};
test_output[3459] = '{32'h42c0cb48};
/*############ DEBUG ############
test_input[27672:27679] = '{-21.6780867042, 14.8391276763, -54.4855223491, -18.0582966643, -80.7052790342, 49.6281767387, 74.7189443718, -33.8281298821};
test_label[3459] = '{-21.6780867042};
test_output[3459] = '{96.397031076};
############ END DEBUG ############*/
test_input[27680:27687] = '{32'h428dce9f, 32'h4214c3d2, 32'h426fb8a7, 32'hc20648bb, 32'hc2aa938e, 32'h40151920, 32'hc22e8fd8, 32'h41d17999};
test_label[3460] = '{32'hc2aa938e};
test_output[3460] = '{32'h431c3117};
/*############ DEBUG ############
test_input[27680:27687] = '{70.903553288, 37.191230046, 59.9303233468, -33.5710266233, -85.2881929851, 2.32965847281, -43.6404723109, 26.1843730368};
test_label[3460] = '{-85.2881929851};
test_output[3460] = '{156.191763428};
############ END DEBUG ############*/
test_input[27688:27695] = '{32'h426a3c7d, 32'hc294677f, 32'h424d86bd, 32'h4202a3a1, 32'hc2b65764, 32'h40bb0e87, 32'hc2581729, 32'hc2bfcef1};
test_label[3461] = '{32'h426a3c7d};
test_output[3461] = '{32'h3a48179a};
/*############ DEBUG ############
test_input[27688:27695] = '{58.5590694381, -74.2021371639, 51.3815801143, 32.6597952903, -91.1706860773, 5.84552314287, -54.0226169556, -95.9041860363};
test_label[3461] = '{58.5590694381};
test_output[3461] = '{0.000763291170889};
############ END DEBUG ############*/
test_input[27696:27703] = '{32'h42bf763d, 32'hc2a35929, 32'hc212dcfe, 32'hc2c5f048, 32'hc1ba2478, 32'hc27cdfe3, 32'hc2870697, 32'h426b3fa0};
test_label[3462] = '{32'hc27cdfe3};
test_output[3462] = '{32'h431ef317};
/*############ DEBUG ############
test_input[27696:27703] = '{95.7309379243, -81.6741397377, -36.7158137541, -98.9693011761, -23.2678060575, -63.2186377211, -67.5128732604, 58.8121350679};
test_label[3462] = '{-63.2186377211};
test_output[3462] = '{158.949575645};
############ END DEBUG ############*/
test_input[27704:27711] = '{32'hc2afcb62, 32'h40b23ae9, 32'hbe4a0e76, 32'hc28736b4, 32'hc1c09f97, 32'hc117b24c, 32'h42b0b9fd, 32'h42840529};
test_label[3463] = '{32'hc2afcb62};
test_output[3463] = '{32'h433042b0};
/*############ DEBUG ############
test_input[27704:27711] = '{-87.8972350822, 5.56969130117, -0.197320784143, -67.6068423505, -24.0779239594, -9.48102964386, 88.3632573556, 66.0100793082};
test_label[3463] = '{-87.8972350822};
test_output[3463] = '{176.260492438};
############ END DEBUG ############*/
test_input[27712:27719] = '{32'h42b8e74e, 32'hc249e2e7, 32'hc23a5878, 32'hc2b916c9, 32'h42bd52c8, 32'hc2977178, 32'hc144247c, 32'hc09a2ec0};
test_label[3464] = '{32'hc144247c};
test_output[3464] = '{32'h42d60ca4};
/*############ DEBUG ############
test_input[27712:27719] = '{92.4517647603, -50.4715856975, -46.586395273, -92.5445048955, 94.6616803148, -75.7216193783, -12.2589077902, -4.81820681442};
test_label[3464] = '{-12.2589077902};
test_output[3464] = '{107.024686746};
############ END DEBUG ############*/
test_input[27720:27727] = '{32'h42c22a45, 32'h428bb6a0, 32'hc285df32, 32'hc18201a3, 32'hc233f2aa, 32'hbf046f62, 32'h42c56435, 32'h41c90354};
test_label[3465] = '{32'h42c22a45};
test_output[3465] = '{32'h3fe5be10};
/*############ DEBUG ############
test_input[27720:27727] = '{97.0825567187, 69.8566874112, -66.935928858, -16.2507996013, -44.9869783445, -0.517324541951, 98.6957174206, 25.1266247406};
test_label[3465] = '{97.0825567187};
test_output[3465] = '{1.79486275543};
############ END DEBUG ############*/
test_input[27728:27735] = '{32'h420591c3, 32'h42bc370f, 32'h42897c8e, 32'h4247d00a, 32'h4228e517, 32'hc2c071b0, 32'h41b925f4, 32'h42a1da78};
test_label[3466] = '{32'h4228e517};
test_output[3466] = '{32'h424f8907};
/*############ DEBUG ############
test_input[27728:27735] = '{33.3923455098, 94.1075353161, 68.7432715177, 49.9531642895, 42.2237196089, -96.2220440069, 23.143531454, 80.9266954505};
test_label[3466] = '{42.2237196089};
test_output[3466] = '{51.8838175936};
############ END DEBUG ############*/
test_input[27736:27743] = '{32'hc2b403db, 32'hc29cdc2c, 32'hc293684d, 32'h42a25dfa, 32'h42833abf, 32'h422c451d, 32'h415241c4, 32'hc1b67c3c};
test_label[3467] = '{32'hc29cdc2c};
test_output[3467] = '{32'h431f9d13};
/*############ DEBUG ############
test_input[27736:27743] = '{-90.0075313474, -78.4300195634, -73.7037099983, 81.1835506086, 65.6147407311, 43.0674946052, 13.1410564086, -22.8106618192};
test_label[3467] = '{-78.4300195634};
test_output[3467] = '{159.613570345};
############ END DEBUG ############*/
test_input[27744:27751] = '{32'h4282e64e, 32'hc1c6b261, 32'h41ee1e74, 32'hc28f42e7, 32'hc2216afa, 32'h42abc7b5, 32'h424327d1, 32'h4061bbe2};
test_label[3468] = '{32'h42abc7b5};
test_output[3468] = '{32'h30b6669f};
/*############ DEBUG ############
test_input[27744:27751] = '{65.4498138215, -24.8370982434, 29.7648697286, -71.6306693953, -40.3544698864, 85.8900527315, 48.7888820199, 3.52709253095};
test_label[3468] = '{85.8900527315};
test_output[3468] = '{1.32714095357e-09};
############ END DEBUG ############*/
test_input[27752:27759] = '{32'hc1e7aa43, 32'hc253a041, 32'hc13cb4af, 32'h4279e459, 32'h4176ff1a, 32'hc20d1746, 32'h428b0b8d, 32'h424dd5e2};
test_label[3469] = '{32'hc20d1746};
test_output[3469] = '{32'h42d197a1};
/*############ DEBUG ############
test_input[27752:27759] = '{-28.958136225, -52.9064997016, -11.7941118869, 62.4729942725, 15.4372803489, -35.2727271846, 69.5225582717, 51.4588691235};
test_label[3469] = '{-35.2727271846};
test_output[3469] = '{104.796152881};
############ END DEBUG ############*/
test_input[27760:27767] = '{32'hc2c2a936, 32'h42c71159, 32'hc071d346, 32'h428b6a0f, 32'h42a3225b, 32'hc2ad8c0c, 32'hc1de6478, 32'hc24ea8f9};
test_label[3470] = '{32'h428b6a0f};
test_output[3470] = '{32'h41ee9d2a};
/*############ DEBUG ############
test_input[27760:27767] = '{-97.3304921675, 99.5338840543, -3.77852003887, 69.7071435349, 81.5671000736, -86.7735325712, -27.799056736, -51.6650116205};
test_label[3470] = '{69.7071435349};
test_output[3470] = '{29.8267405352};
############ END DEBUG ############*/
test_input[27768:27775] = '{32'hc29ad11e, 32'hc2c510a6, 32'hc2bafc19, 32'h40bf32ab, 32'h429fb391, 32'h42ab6e56, 32'h429b8fc2, 32'hc2948a7b};
test_label[3471] = '{32'hc29ad11e};
test_output[3471] = '{32'h4323208b};
/*############ DEBUG ############
test_input[27768:27775] = '{-77.4084285462, -98.5325194819, -93.492377795, 5.97493493527, 79.8507153921, 85.7154994855, 77.7807736726, -74.2704699999};
test_label[3471] = '{-77.4084285462};
test_output[3471] = '{163.127118662};
############ END DEBUG ############*/
test_input[27776:27783] = '{32'hc2b0b5e6, 32'h42400c2a, 32'hc218a87f, 32'hc101f181, 32'h420cb557, 32'h4238d6e3, 32'h42b255bb, 32'h41c5bc89};
test_label[3472] = '{32'h420cb557};
test_output[3472] = '{32'h4257f61e};
/*############ DEBUG ############
test_input[27776:27783] = '{-88.3552728299, 48.0118792223, -38.1645475072, -8.12146059887, 35.1770901638, 46.2098487748, 89.1674389626, 24.7170589505};
test_label[3472] = '{35.1770901638};
test_output[3472] = '{53.9903487988};
############ END DEBUG ############*/
test_input[27784:27791] = '{32'h428807c5, 32'hc2ade3ca, 32'hc19d0e71, 32'h42b22c01, 32'h42865a87, 32'hc2209ea7, 32'hc2c48196, 32'h423c666c};
test_label[3473] = '{32'h42b22c01};
test_output[3473] = '{32'h308b142f};
/*############ DEBUG ############
test_input[27784:27791] = '{68.0151740321, -86.9449019166, -19.6320521257, 89.0859424231, 67.1768110133, -40.1549344942, -98.2530946371, 47.1000203438};
test_label[3473] = '{89.0859424231};
test_output[3473] = '{1.01193176112e-09};
############ END DEBUG ############*/
test_input[27792:27799] = '{32'hc2ba79b7, 32'hc2ab0f47, 32'hc2a49c08, 32'h41d3249b, 32'hc2167f85, 32'hc1cf0f78, 32'h41aad602, 32'h406ce9d7};
test_label[3474] = '{32'h41d3249b};
test_output[3474] = '{32'h3bd3ca54};
/*############ DEBUG ############
test_input[27792:27799] = '{-93.2377218527, -85.5298368656, -82.3047464489, 26.3928728758, -37.6245306342, -25.8825531094, 21.3544954161, 3.70177247585};
test_label[3474] = '{26.3928728758};
test_output[3474] = '{0.00646332852042};
############ END DEBUG ############*/
test_input[27800:27807] = '{32'h4199558c, 32'hc2bc24e8, 32'hc11f5fb6, 32'h423d5e30, 32'hc23d987f, 32'hc1c012de, 32'h42562388, 32'h427b2649};
test_label[3475] = '{32'hc11f5fb6};
test_output[3475] = '{32'h42917f28};
/*############ DEBUG ############
test_input[27800:27807] = '{19.1667711399, -94.0720835134, -9.96086691409, 47.3419811602, -47.3989216154, -24.0092123625, 53.5346975817, 62.7873872759};
test_label[3475] = '{-9.96086691409};
test_output[3475] = '{72.7483502348};
############ END DEBUG ############*/
test_input[27808:27815] = '{32'hc131ebec, 32'hc0d1aeb2, 32'h429ffae2, 32'hc2bad7f0, 32'hc19348ee, 32'h42c545b6, 32'h4103ab54, 32'h4218f23d};
test_label[3476] = '{32'h4218f23d};
test_output[3476] = '{32'h4271992f};
/*############ DEBUG ############
test_input[27808:27815] = '{-11.120097936, -6.55257504683, 79.9900031522, -93.4217533664, -18.4106097469, 98.6361546861, 8.22932824996, 38.2365615563};
test_label[3476] = '{38.2365615563};
test_output[3476] = '{60.3995931378};
############ END DEBUG ############*/
test_input[27816:27823] = '{32'hc2792243, 32'hc2b8b55e, 32'hc219906e, 32'hc20d042b, 32'h421cdf7e, 32'hc20325b3, 32'hc2b1636c, 32'hc2a3a8a2};
test_label[3477] = '{32'hc2792243};
test_output[3477] = '{32'h42cb00e1};
/*############ DEBUG ############
test_input[27816:27823] = '{-62.2834595617, -92.3542359456, -38.3910442095, -35.2540692115, 39.2182554878, -32.7868147602, -88.6941824937, -81.8293600244};
test_label[3477] = '{-62.2834595617};
test_output[3477] = '{101.501715049};
############ END DEBUG ############*/
test_input[27824:27831] = '{32'hc297f64a, 32'hc2815d4d, 32'h41b77804, 32'hc21b566d, 32'h41e2b309, 32'h42c62f79, 32'hc264e7fe, 32'hc219287e};
test_label[3478] = '{32'h41b77804};
test_output[3478] = '{32'h42985178};
/*############ DEBUG ############
test_input[27824:27831] = '{-75.9810323074, -64.6822314636, 22.9336010789, -38.8343991422, 28.337419179, 99.0927202712, -57.2265545418, -38.289541601};
test_label[3478] = '{22.9336010789};
test_output[3478] = '{76.1591191923};
############ END DEBUG ############*/
test_input[27832:27839] = '{32'h41e4beb1, 32'h42097560, 32'hc2c3b54c, 32'hc224b67a, 32'hc2c6e6b1, 32'hc2732756, 32'h41c7b4f1, 32'h417ae27d};
test_label[3479] = '{32'h42097560};
test_output[3479] = '{32'h3b513a61};
/*############ DEBUG ############
test_input[27832:27839] = '{28.5931101627, 34.3646228964, -97.8540962178, -41.1782006507, -99.450571703, -60.788413684, 24.963351002, 15.6802946196};
test_label[3479] = '{34.3646228964};
test_output[3479] = '{0.00319256664975};
############ END DEBUG ############*/
test_input[27840:27847] = '{32'hc2a7ea08, 32'h4227a0d8, 32'h42ae9df1, 32'h42c4a5ae, 32'hc2b0e238, 32'h42062ede, 32'h41b0b8ca, 32'h42b4cf25};
test_label[3480] = '{32'h42062ede};
test_output[3480] = '{32'h42818e71};
/*############ DEBUG ############
test_input[27840:27847] = '{-83.9570908073, 41.907075055, 87.3084767765, 98.3235928179, -88.4418342197, 33.5457700876, 22.0902288291, 90.4045822533};
test_label[3480] = '{33.5457700876};
test_output[3480] = '{64.7782028712};
############ END DEBUG ############*/
test_input[27848:27855] = '{32'h4285177e, 32'h4278b8ec, 32'hc230ed8c, 32'h41b3ef3e, 32'hc2bf224b, 32'hc1af0dfb, 32'hc200b92e, 32'hc2a7220f};
test_label[3481] = '{32'hc200b92e};
test_output[3481] = '{32'h42c57a8d};
/*############ DEBUG ############
test_input[27848:27855] = '{66.545886104, 62.1805867191, -44.231978857, 22.4918167644, -95.5669820129, -21.8818257509, -32.1808403229, -83.5665226111};
test_label[3481] = '{-32.1808403229};
test_output[3481] = '{98.7393571713};
############ END DEBUG ############*/
test_input[27856:27863] = '{32'hc2bb565b, 32'h412502fc, 32'h41a02a61, 32'h41cf0087, 32'hc27ed413, 32'hc1c95849, 32'h42480987, 32'h425fce07};
test_label[3482] = '{32'hc2bb565b};
test_output[3482] = '{32'h43159f5b};
/*############ DEBUG ############
test_input[27856:27863] = '{-93.6686615987, 10.3132287926, 20.0206931409, 25.8752567949, -63.7071024696, -25.1681076448, 50.0093048231, 55.9511987766};
test_label[3482] = '{-93.6686615987};
test_output[3482] = '{149.62248398};
############ END DEBUG ############*/
test_input[27864:27871] = '{32'hc2b61bf7, 32'h3f14a4a6, 32'h421b85a3, 32'h42bf2e61, 32'h4180b2ee, 32'h42bf0150, 32'hc2bbbc25, 32'h425d70ad};
test_label[3483] = '{32'h421b85a3};
test_output[3483] = '{32'h426570d5};
/*############ DEBUG ############
test_input[27864:27871] = '{-91.054619911, 0.58063731248, 38.880503109, 95.5905867558, 16.0873679882, 95.5025659243, -93.8674712067, 55.360036644};
test_label[3483] = '{38.880503109};
test_output[3483] = '{57.3601885575};
############ END DEBUG ############*/
test_input[27872:27879] = '{32'hc14e03ba, 32'h4208233a, 32'h42be2cf5, 32'h402fd52b, 32'hc2a47a65, 32'h42497d44, 32'h42aaec95, 32'hc28d128d};
test_label[3484] = '{32'hc28d128d};
test_output[3484] = '{32'h43259fc5};
/*############ DEBUG ############
test_input[27872:27879] = '{-12.8759097389, 34.034401917, 95.0878032597, 2.74738566837, -82.2390496726, 50.3723278159, 85.4620751044, -70.5362349043};
test_label[3484] = '{-70.5362349043};
test_output[3484] = '{165.62410417};
############ END DEBUG ############*/
test_input[27880:27887] = '{32'h4248cd2f, 32'hc2667150, 32'h42b9a7bc, 32'h428d819b, 32'hc1bfbbdc, 32'h42b8ecb8, 32'h42c14d08, 32'hc21c067f};
test_label[3485] = '{32'hc1bfbbdc};
test_output[3485] = '{32'h42f14e9f};
/*############ DEBUG ############
test_input[27880:27887] = '{50.2003755996, -57.6106573449, 92.8276031093, 70.7531321653, -23.9667277452, 92.4623432673, 96.6504545497, -39.0063453805};
test_label[3485] = '{-23.9667277452};
test_output[3485] = '{120.653553069};
############ END DEBUG ############*/
test_input[27888:27895] = '{32'h42099f79, 32'h41eacee6, 32'h407a53c6, 32'h41fc8bc1, 32'h41b43c1f, 32'h418ba03d, 32'hc24bedcd, 32'hc0504794};
test_label[3486] = '{32'h418ba03d};
test_output[3486] = '{32'h41881f99};
/*############ DEBUG ############
test_input[27888:27895] = '{34.4057349435, 29.3510245545, 3.91136323213, 31.5682388643, 22.5293564768, 17.4532414927, -50.9822268836, -3.25436880023};
test_label[3486] = '{17.4532414927};
test_output[3486] = '{17.0154291437};
############ END DEBUG ############*/
test_input[27896:27903] = '{32'hc205f6f1, 32'h4188b470, 32'h419c7331, 32'h42aac3dd, 32'h401e2696, 32'hc18e4701, 32'hc1f11841, 32'h41fc3fc1};
test_label[3487] = '{32'hc18e4701};
test_output[3487] = '{32'h42ce559d};
/*############ DEBUG ############
test_input[27896:27903] = '{-33.4911552767, 17.0881042067, 19.5562459918, 85.3825433297, 2.47110499092, -17.784669693, -30.136842131, 31.5311302313};
test_label[3487] = '{-17.784669693};
test_output[3487] = '{103.167213023};
############ END DEBUG ############*/
test_input[27904:27911] = '{32'hc296812a, 32'hc269e142, 32'h42b3c8a0, 32'h4260bcdf, 32'hc23417b6, 32'hc280447a, 32'h4280e926, 32'h429b7b08};
test_label[3488] = '{32'hc269e142};
test_output[3488] = '{32'h43145ca1};
/*############ DEBUG ############
test_input[27904:27911] = '{-75.252272022, -58.4699794104, 89.8918474192, 56.1844451822, -45.0231552815, -64.1337462648, 64.4553701288, 77.7402956203};
test_label[3488] = '{-58.4699794104};
test_output[3488] = '{148.36183211};
############ END DEBUG ############*/
test_input[27912:27919] = '{32'h429078ae, 32'hc24c5ea4, 32'h40e00751, 32'h41c90158, 32'hc242c4bb, 32'hc2a61105, 32'h4282ed10, 32'h42b7f0ca};
test_label[3489] = '{32'h429078ae};
test_output[3489] = '{32'h419de06f};
/*############ DEBUG ############
test_input[27912:27919] = '{72.2357034512, -51.0924219742, 7.00089293526, 25.1256563822, -48.6921191343, -83.0332414116, 65.4630101563, 91.9702895593};
test_label[3489] = '{72.2357034512};
test_output[3489] = '{19.7345861108};
############ END DEBUG ############*/
test_input[27920:27927] = '{32'h40d30b2a, 32'hc24f6b4a, 32'h426a1703, 32'hc2bef180, 32'h420cf92c, 32'h41593003, 32'h42a8315f, 32'hc2b78563};
test_label[3490] = '{32'h40d30b2a};
test_output[3490] = '{32'h429b00ac};
/*############ DEBUG ############
test_input[27920:27927] = '{6.59511294053, -51.8547734799, 58.5224721301, -95.4716776771, 35.2433323045, 13.5742212872, 84.0964282378, -91.760517453};
test_label[3490] = '{6.59511294053};
test_output[3490] = '{77.5013152973};
############ END DEBUG ############*/
test_input[27928:27935] = '{32'h4058340c, 32'h421e5921, 32'hc2ab4c7c, 32'h429e6ad8, 32'h42c25445, 32'hc2375226, 32'h42b53d81, 32'hc236b211};
test_label[3491] = '{32'h429e6ad8};
test_output[3491] = '{32'h418fa8a6};
/*############ DEBUG ############
test_input[27928:27935] = '{3.37817674564, 39.5870399589, -85.6493803867, 79.2086771355, 97.1645871777, -45.8302246371, 90.6201221467, -45.6738945511};
test_label[3491] = '{79.2086771355};
test_output[3491] = '{17.9573470782};
############ END DEBUG ############*/
test_input[27936:27943] = '{32'hc2c07513, 32'h42c15e0e, 32'h428feb99, 32'hc2a3dc1d, 32'hc2b7895a, 32'h428fa5b1, 32'h411245b5, 32'hc2b91e98};
test_label[3492] = '{32'hc2b7895a};
test_output[3492] = '{32'h433c73b4};
/*############ DEBUG ############
test_input[27936:27943] = '{-96.2286628868, 96.6837001916, 71.9601547531, -81.9299090005, -91.7682641105, 71.8236194297, 9.14201814333, -92.5597562318};
test_label[3492] = '{-91.7682641105};
test_output[3492] = '{188.451964302};
############ END DEBUG ############*/
test_input[27944:27951] = '{32'hc2c6865b, 32'h42c52704, 32'h427ac002, 32'h429c3372, 32'h42a33480, 32'h423b747b, 32'h4084b8b0, 32'h42397532};
test_label[3493] = '{32'h423b747b};
test_output[3493] = '{32'h424ed98c};
/*############ DEBUG ############
test_input[27944:27951] = '{-99.2624099454, 98.5761990224, 62.6875074169, 78.100479956, 81.6025415544, 46.8637516586, 4.14754508591, 46.364448185};
test_label[3493] = '{46.8637516586};
test_output[3493] = '{51.7124474076};
############ END DEBUG ############*/
test_input[27952:27959] = '{32'hc1fc5356, 32'hc0b4bd68, 32'hc29f599f, 32'h42299c2a, 32'h4271d76d, 32'h422eb6e7, 32'h42872695, 32'hc24c8c3a};
test_label[3494] = '{32'h42299c2a};
test_output[3494] = '{32'h41c963ab};
/*############ DEBUG ############
test_input[27952:27959] = '{-31.5406920087, -5.64812111753, -79.6750379696, 42.4025031077, 60.4603770265, 43.6786168371, 67.5753567024, -51.1369401632};
test_label[3494] = '{42.4025031077};
test_output[3494] = '{25.1736661018};
############ END DEBUG ############*/
test_input[27960:27967] = '{32'hc2382424, 32'h3f91338a, 32'h423a445b, 32'hc11b3fc2, 32'hc2a353b2, 32'hc18011f4, 32'hc23c6831, 32'h4229f3f5};
test_label[3495] = '{32'hc23c6831};
test_output[3495] = '{32'h42bb5edf};
/*############ DEBUG ############
test_input[27960:27967] = '{-46.0352934687, 1.13438536954, 46.5667527132, -9.70306610063, -81.6634702108, -16.0087668157, -47.1017502778, 42.488239405};
test_label[3495] = '{-47.1017502778};
test_output[3495] = '{93.6852938527};
############ END DEBUG ############*/
test_input[27968:27975] = '{32'hc2c07b98, 32'h428f71eb, 32'hc28e6b3b, 32'hc29dd601, 32'h41cd0401, 32'hc15d5ad9, 32'h423f5b82, 32'hc2be9fce};
test_label[3496] = '{32'h41cd0401};
test_output[3496] = '{32'h423861d5};
/*############ DEBUG ############
test_input[27968:27975] = '{-96.2413958636, 71.7224934874, -71.2094348625, -78.91797864, 25.6269547956, -13.8346799062, 47.8393649471, -95.3121215612};
test_label[3496] = '{25.6269547956};
test_output[3496] = '{46.0955386919};
############ END DEBUG ############*/
test_input[27976:27983] = '{32'hc10cb044, 32'hc2b51ef6, 32'h41f796e9, 32'h427f8fe6, 32'h41464453, 32'h41e0c711, 32'h4285d905, 32'hc2a8fa01};
test_label[3497] = '{32'h4285d905};
test_output[3497] = '{32'h3d40a395};
/*############ DEBUG ############
test_input[27976:27983] = '{-8.79303361825, -90.5604734493, 30.9486860202, 63.8905258301, 12.391680608, 28.0972008899, 66.9238663885, -84.4882867267};
test_label[3497] = '{66.9238663885};
test_output[3497] = '{0.0470310046148};
############ END DEBUG ############*/
test_input[27984:27991] = '{32'h42818dac, 32'h420611f6, 32'h42791a19, 32'h42c5ddf8, 32'hc29f7c2f, 32'hc222f391, 32'hc082aad9, 32'h42ba332b};
test_label[3498] = '{32'hc29f7c2f};
test_output[3498] = '{32'h4332add3};
/*############ DEBUG ############
test_input[27984:27991] = '{64.7767041172, 33.5175412251, 62.2754858118, 98.9335344545, -79.7425456437, -40.7378590536, -4.08335556303, 93.0999364066};
test_label[3498] = '{-79.7425456437};
test_output[3498] = '{178.679003346};
############ END DEBUG ############*/
test_input[27992:27999] = '{32'h4261cccb, 32'h41af84ae, 32'h41c7c203, 32'h42969652, 32'hc20bdb80, 32'h41941266, 32'h4250dae3, 32'hc1d40be6};
test_label[3499] = '{32'hc1d40be6};
test_output[3499] = '{32'h42cb994c};
/*############ DEBUG ############
test_input[27992:27999] = '{56.4499940191, 21.9397853783, 24.9697328615, 75.2935979796, -34.9643553143, 18.5089835871, 52.2137552107, -26.5058097638};
test_label[3499] = '{-26.5058097638};
test_output[3499] = '{101.79940775};
############ END DEBUG ############*/
test_input[28000:28007] = '{32'h422153f5, 32'hc204b81e, 32'h42c38e89, 32'h420c2a7c, 32'h42aa01a3, 32'h4166f949, 32'h41f77bf6, 32'h4238c38c};
test_label[3500] = '{32'h42aa01a3};
test_output[3500] = '{32'h414c6737};
/*############ DEBUG ############
test_input[28000:28007] = '{40.3319910054, -33.1798019876, 97.7783924128, 35.041488905, 85.003196304, 14.4358610227, 30.9355268515, 46.1909628353};
test_label[3500] = '{85.003196304};
test_output[3500] = '{12.7751989389};
############ END DEBUG ############*/
test_input[28008:28015] = '{32'h4134c98f, 32'h423ecfdb, 32'hc0b15509, 32'hbf0f1ada, 32'hc2808b27, 32'h428051af, 32'hc2814412, 32'h42aa14dc};
test_label[3501] = '{32'h428051af};
test_output[3501] = '{32'h41a70cb6};
/*############ DEBUG ############
test_input[28008:28015] = '{11.2992084455, 47.7029835121, -5.54163041055, -0.559003448238, -64.271784037, 64.159535994, -64.6329512155, 85.0407430412};
test_label[3501] = '{64.159535994};
test_output[3501] = '{20.881207048};
############ END DEBUG ############*/
test_input[28016:28023] = '{32'hc2bbe874, 32'hc1237708, 32'h425e7968, 32'hc1658d30, 32'h423d62e4, 32'hc21f1a56, 32'h420e39cf, 32'hc1750f64};
test_label[3502] = '{32'h420e39cf};
test_output[3502] = '{32'h41a07fb7};
/*############ DEBUG ############
test_input[28016:28023] = '{-93.9540100641, -10.2165607264, 55.6185592094, -14.3469693188, 47.3465741792, -39.7757200497, 35.5564542272, -15.3162570116};
test_label[3502] = '{35.5564542272};
test_output[3502] = '{20.0623605289};
############ END DEBUG ############*/
test_input[28024:28031] = '{32'hc1ea6ffd, 32'hc2b4b0a9, 32'h428d1a52, 32'hc1945335, 32'h428c4d3d, 32'h42b18e9a, 32'hc2b3f39f, 32'hc23a11a4};
test_label[3503] = '{32'h42b18e9a};
test_output[3503] = '{32'h32ae15ab};
/*############ DEBUG ############
test_input[28024:28031] = '{-29.3046819542, -90.3450386993, 70.5514062178, -18.5406288698, 70.1508568103, 88.7785163028, -89.9758255022, -46.5172254589};
test_label[3503] = '{88.7785163028};
test_output[3503] = '{2.02661203208e-08};
############ END DEBUG ############*/
test_input[28032:28039] = '{32'hc2897991, 32'hc2ac3c9c, 32'h4218db3c, 32'h41a30b7b, 32'h4249cc6f, 32'h413b2e2a, 32'h42bc8655, 32'hc2b44616};
test_label[3504] = '{32'hc2b44616};
test_output[3504] = '{32'h43386636};
/*############ DEBUG ############
test_input[28032:28039] = '{-68.7374355912, -86.1183806998, 38.2140963577, 20.3806053434, 50.4496412423, 11.6987702789, 94.2623651009, -90.1368892681};
test_label[3504] = '{-90.1368892681};
test_output[3504] = '{184.399254369};
############ END DEBUG ############*/
test_input[28040:28047] = '{32'hc2521c33, 32'hc287cf1d, 32'hc29d270e, 32'h40a3a8b2, 32'hc2512c6c, 32'h42c31c5a, 32'h429aad73, 32'h424b48d5};
test_label[3505] = '{32'h42c31c5a};
test_output[3505] = '{32'h30e41d24};
/*############ DEBUG ############
test_input[28040:28047] = '{-52.5275380633, -67.9045151715, -78.5762776098, 5.11434246927, -52.2933826316, 97.5553717523, 77.3387708234, 50.8211266764};
test_label[3505] = '{97.5553717523};
test_output[3505] = '{1.65974656379e-09};
############ END DEBUG ############*/
test_input[28048:28055] = '{32'hc22b87f8, 32'h411263d9, 32'hc2b350bb, 32'h41e5a454, 32'hc214ba11, 32'h41710bee, 32'h4276b5e3, 32'hc176b58e};
test_label[3506] = '{32'h41e5a454};
test_output[3506] = '{32'h4203e3b9};
/*############ DEBUG ############
test_input[28048:28055] = '{-42.8827825034, 9.14937718082, -89.6576750438, 28.7052388833, -37.1817064337, 15.0654122854, 61.677623517, -15.4193248122};
test_label[3506] = '{28.7052388833};
test_output[3506] = '{32.9723846338};
############ END DEBUG ############*/
test_input[28056:28063] = '{32'hc1b652e2, 32'h4293a904, 32'h40d1137d, 32'hc294f27a, 32'h42a282a2, 32'h42b8474d, 32'hc1bc0031, 32'hc2be188f};
test_label[3507] = '{32'hc2be188f};
test_output[3507] = '{32'h433b2fef};
/*############ DEBUG ############
test_input[28056:28063] = '{-22.7904709358, 73.8301048638, 6.53362872439, -74.473587694, 81.2551449332, 92.1392623306, -23.5000930237, -95.0479635732};
test_label[3507] = '{-95.0479635732};
test_output[3507] = '{187.187244669};
############ END DEBUG ############*/
test_input[28064:28071] = '{32'hc2bb6e58, 32'h42351fb8, 32'h423fca13, 32'hc28421b6, 32'h4284ed22, 32'h420725fb, 32'hc181ce8f, 32'h4018e6bd};
test_label[3508] = '{32'hc28421b6};
test_output[3508] = '{32'h4304876c};
/*############ DEBUG ############
test_input[28064:28071] = '{-93.7155130469, 45.2809766457, 47.9473377689, -66.0658445969, 66.4631468037, 33.7870891789, -16.2258584644, 2.38908314589};
test_label[3508] = '{-66.0658445969};
test_output[3508] = '{132.52899141};
############ END DEBUG ############*/
test_input[28072:28079] = '{32'hc1cf5acf, 32'hc2a91f79, 32'hc1f447bd, 32'hc1ace937, 32'hc1883f0f, 32'h41fd733f, 32'h42a9deb1, 32'h4190c177};
test_label[3509] = '{32'hc1883f0f};
test_output[3509] = '{32'h42cbee75};
/*############ DEBUG ############
test_input[28072:28079] = '{-25.9193409173, -84.5614697031, -30.535029201, -21.6138749991, -17.0307903189, 31.6812730371, 84.9349435046, 18.0944644648};
test_label[3509] = '{-17.0307903189};
test_output[3509] = '{101.965733823};
############ END DEBUG ############*/
test_input[28080:28087] = '{32'hc2964319, 32'h40ffb01b, 32'h42769802, 32'h41c52a38, 32'h41ac20b1, 32'hc27854d5, 32'h42b4cfc0, 32'hc0f64db3};
test_label[3510] = '{32'hc27854d5};
test_output[3510] = '{32'h43187d16};
/*############ DEBUG ############
test_input[28080:28087] = '{-75.1310463194, 7.9902473119, 61.6484460092, 24.6456144718, 21.5159632885, -62.0828454506, 90.4057653293, -7.69698490883};
test_label[3510] = '{-62.0828454506};
test_output[3510] = '{152.48861078};
############ END DEBUG ############*/
test_input[28088:28095] = '{32'hc1e92225, 32'h42212a9f, 32'h421915c5, 32'h41ea882e, 32'h3fe917c8, 32'h4264d6d9, 32'h428068ce, 32'h42781188};
test_label[3511] = '{32'hc1e92225};
test_output[3511] = '{32'h42bae834};
/*############ DEBUG ############
test_input[28088:28095] = '{-29.1416727657, 40.2916221905, 38.2712602572, 29.3164945149, 1.82103823539, 57.2098110032, 64.2046939332, 62.017119765};
test_label[3511] = '{-29.1416727657};
test_output[3511] = '{93.4535202227};
############ END DEBUG ############*/
test_input[28096:28103] = '{32'hc24f69b7, 32'h3e1cd74d, 32'h42c75663, 32'h422187f8, 32'h4292a238, 32'hc2a48959, 32'hc268683a, 32'h4082f687};
test_label[3512] = '{32'h4082f687};
test_output[3512] = '{32'h42bf26fb};
/*############ DEBUG ############
test_input[28096:28103] = '{-51.8532364375, 0.15316505559, 99.6687265466, 40.3827811906, 73.3168334918, -82.2682551098, -58.1017841945, 4.09259377106};
test_label[3512] = '{4.09259377106};
test_output[3512] = '{95.5761327755};
############ END DEBUG ############*/
test_input[28104:28111] = '{32'h41e17078, 32'h41fb66cf, 32'hc273227f, 32'h41493cbe, 32'hc20f0f32, 32'h429a4a0c, 32'hc2c162cb, 32'hc2c43dc7};
test_label[3513] = '{32'hc2c162cb};
test_output[3513] = '{32'h432dd66c};
/*############ DEBUG ############
test_input[28104:28111] = '{28.1799154859, 31.4251999158, -60.7836887855, 12.5773299469, -35.7648375067, 77.1446259608, -96.6929521949, -98.120657136};
test_label[3513] = '{-96.6929521949};
test_output[3513] = '{173.837578156};
############ END DEBUG ############*/
test_input[28112:28119] = '{32'hc2854e67, 32'h4203ceff, 32'hc2c189ff, 32'h4105a7fb, 32'h42832e18, 32'hc2adf566, 32'h42b7487d, 32'h42b55242};
test_label[3514] = '{32'hc2adf566};
test_output[3514] = '{32'h4332f076};
/*############ DEBUG ############
test_input[28112:28119] = '{-66.6531325207, 32.9521431166, -96.7695272214, 8.35351047406, 65.5900256038, -86.9792905954, 91.6415775209, 90.6606603537};
test_label[3514] = '{-86.9792905954};
test_output[3514] = '{178.939297872};
############ END DEBUG ############*/
test_input[28120:28127] = '{32'h42c66f0a, 32'h42a01d4f, 32'hc2b8fb46, 32'hc2abb80d, 32'hc211a9f1, 32'hc2ae49d6, 32'hc1427eb5, 32'h41f8792e};
test_label[3515] = '{32'hc1427eb5};
test_output[3515] = '{32'h42debee1};
/*############ DEBUG ############
test_input[28120:28127] = '{99.2168734651, 80.0572432274, -92.4907698128, -85.8594764782, -36.4159582122, -87.1442141051, -12.1559343814, 31.0591699395};
test_label[3515] = '{-12.1559343814};
test_output[3515] = '{111.372807851};
############ END DEBUG ############*/
test_input[28128:28135] = '{32'h4249100f, 32'h42ae8c2e, 32'hc24ca782, 32'hc1d19b0a, 32'hc19784fe, 32'hc15c1ff3, 32'h419f4204, 32'h418c19be};
test_label[3516] = '{32'h418c19be};
test_output[3516] = '{32'h428b85bf};
/*############ DEBUG ############
test_input[28128:28135] = '{50.2656821566, 87.2737894274, -51.1635810729, -26.2007031438, -18.9399384108, -13.7578002139, 19.9072336552, 17.5125699012};
test_label[3516] = '{17.5125699012};
test_output[3516] = '{69.7612195261};
############ END DEBUG ############*/
test_input[28136:28143] = '{32'hc1c3b699, 32'hc25ad553, 32'h423b3b24, 32'hc2700761, 32'hc2aedb30, 32'hc221fc8d, 32'h429c6ad7, 32'h425b5a9f};
test_label[3517] = '{32'h429c6ad7};
test_output[3517] = '{32'h2e9be560};
/*############ DEBUG ############
test_input[28136:28143] = '{-24.4641597213, -54.7083240706, 46.8077552879, -60.0072041097, -87.428097095, -40.4966330034, 78.2086697276, 54.8384975794};
test_label[3517] = '{78.2086697276};
test_output[3517] = '{7.089329124e-11};
############ END DEBUG ############*/
test_input[28144:28151] = '{32'hc211a1cf, 32'hc296961e, 32'h41821730, 32'h424ede22, 32'hc286a119, 32'h4108effb, 32'hc291c15d, 32'hc2814b8b};
test_label[3518] = '{32'h424ede22};
test_output[3518] = '{32'h26000000};
/*############ DEBUG ############
test_input[28144:28151] = '{-36.4080155305, -75.2931985416, 16.2613221336, 51.7169264084, -67.3146412541, 8.55858860487, -72.8776601241, -64.6475440971};
test_label[3518] = '{51.7169264084};
test_output[3518] = '{4.4408920985e-16};
############ END DEBUG ############*/
test_input[28152:28159] = '{32'hc25042f4, 32'hc21e6000, 32'hc1651c7b, 32'hc11730ee, 32'h421aabd1, 32'h41b0ed77, 32'hc2b8b6a4, 32'h4297fe1d};
test_label[3519] = '{32'hc21e6000};
test_output[3519] = '{32'h42e72e1d};
/*############ DEBUG ############
test_input[28152:28159] = '{-52.0653832926, -39.5937508246, -14.3194532968, -9.44944605027, 38.6677910675, 22.1159503808, -92.356723254, 75.9963132925};
test_label[3519] = '{-39.5937508246};
test_output[3519] = '{115.590064117};
############ END DEBUG ############*/
test_input[28160:28167] = '{32'h40fbd16b, 32'h41e20699, 32'hc033d771, 32'hc2708d48, 32'h42605d79, 32'h408b16f9, 32'hc2330c75, 32'hc1280dc0};
test_label[3520] = '{32'hc1280dc0};
test_output[3520] = '{32'h42853074};
/*############ DEBUG ############
test_input[28160:28167] = '{7.86931352542, 28.253221862, -2.81002441395, -60.1379684188, 56.091280774, 4.34655423502, -44.7621648969, -10.5033564962};
test_label[3520] = '{-10.5033564962};
test_output[3520] = '{66.5946372702};
############ END DEBUG ############*/
test_input[28168:28175] = '{32'hc164abd0, 32'hbf89c2a2, 32'hc23486d9, 32'hc22bf282, 32'h413d7471, 32'hc2bf12ef, 32'h40d45bab, 32'h419bc7a4};
test_label[3521] = '{32'hbf89c2a2};
test_output[3521] = '{32'h41a464ce};
/*############ DEBUG ############
test_input[28168:28175] = '{-14.2919465995, -1.07625224566, -45.1316866018, -42.9868242184, 11.8409278117, -95.5369778966, 6.6361900452, 19.4724807205};
test_label[3521] = '{-1.07625224566};
test_output[3521] = '{20.5492204181};
############ END DEBUG ############*/
test_input[28176:28183] = '{32'h42b053f1, 32'hc2c45b8b, 32'h4205cb82, 32'hc2ac23a5, 32'hc271fcc0, 32'hc1588188, 32'h405e6e9a, 32'hc2a8ec28};
test_label[3522] = '{32'hc1588188};
test_output[3522] = '{32'h42cb6422};
/*############ DEBUG ############
test_input[28176:28183] = '{88.1639483143, -98.1787940607, 33.4487393808, -86.0696214648, -60.4968244646, -13.5316233987, 3.4755005743, -84.4612421183};
test_label[3522] = '{-13.5316233987};
test_output[3522] = '{101.695571713};
############ END DEBUG ############*/
test_input[28184:28191] = '{32'h42af30a7, 32'h40445f4e, 32'hc284c541, 32'h428f1cf5, 32'h42536219, 32'h41c19ca0, 32'hc2be4de1, 32'h429fe15d};
test_label[3523] = '{32'h428f1cf5};
test_output[3523] = '{32'h41804fc1};
/*############ DEBUG ############
test_input[28184:28191] = '{87.5950237746, 3.06831704246, -66.3852592902, 71.556554775, 52.8457969349, 24.2014761618, -95.1521110232, 79.9401661993};
test_label[3523] = '{71.556554775};
test_output[3523] = '{16.038942733};
############ END DEBUG ############*/
test_input[28192:28199] = '{32'h3f859b7e, 32'hc156cd22, 32'hc2675d48, 32'h42b9039d, 32'h41ddebc1, 32'h41eab7b4, 32'h42a57c37, 32'h41a653d3};
test_label[3524] = '{32'h41a653d3};
test_output[3524] = '{32'h428f6eb0};
/*############ DEBUG ############
test_input[28192:28199] = '{1.04380774699, -13.4250811905, -57.8410934889, 92.5070603339, 27.7401134026, 29.3396996622, 82.742608016, 20.7909301231};
test_label[3524] = '{20.7909301231};
test_output[3524] = '{71.7161876675};
############ END DEBUG ############*/
test_input[28200:28207] = '{32'hc1d5bc5c, 32'hc162344a, 32'h400d2756, 32'h413b4085, 32'hc2870dbd, 32'hc2104606, 32'hc2bbf2a9, 32'h41c0f477};
test_label[3525] = '{32'h41c0f477};
test_output[3525] = '{32'h3687ff64};
/*############ DEBUG ############
test_input[28200:28207] = '{-26.7169727512, -14.1377658359, 2.20552584867, 11.7032517144, -67.5268306857, -36.0683805861, -93.9739450694, 24.1193668903};
test_label[3525] = '{24.1193668903};
test_output[3525] = '{4.05304469401e-06};
############ END DEBUG ############*/
test_input[28208:28215] = '{32'h4196b9d9, 32'h41d81b9a, 32'hc0999d55, 32'hc23ede4c, 32'h42c67772, 32'h41c35c88, 32'h41cb0a78, 32'hc18a1d44};
test_label[3526] = '{32'hc18a1d44};
test_output[3526] = '{32'h42e8fec3};
/*############ DEBUG ############
test_input[28208:28215] = '{18.8407456423, 27.0134782401, -4.80045543896, -47.7170881532, 99.2332927533, 24.4201810323, 25.3801123087, -17.2642898907};
test_label[3526] = '{-17.2642898907};
test_output[3526] = '{116.497582644};
############ END DEBUG ############*/
test_input[28216:28223] = '{32'h42aab4af, 32'h41d308b9, 32'h423c017f, 32'hc12ea5af, 32'h428de276, 32'hc2a15580, 32'h4149b6ad, 32'h422fc366};
test_label[3527] = '{32'h428de276};
test_output[3527] = '{32'h416691cd};
/*############ DEBUG ############
test_input[28216:28223] = '{85.3528995983, 26.3792595671, 47.0014591263, -10.9154496799, 70.9423044764, -80.6669917485, 12.6070990215, 43.9408181012};
test_label[3527] = '{70.9423044764};
test_output[3527] = '{14.4105956734};
############ END DEBUG ############*/
test_input[28224:28231] = '{32'h401173fa, 32'hc2246c50, 32'hc0cad334, 32'h409252c6, 32'h4155979a, 32'h42b8d069, 32'hc2af0048, 32'hc23eee82};
test_label[3528] = '{32'h409252c6};
test_output[3528] = '{32'h42afab3c};
/*############ DEBUG ############
test_input[28224:28231] = '{2.2727037048, -41.1057736063, -6.33828168443, 4.57260404814, 13.3495121814, 92.407047538, -87.5005517923, -47.7329184756};
test_label[3528] = '{4.57260404814};
test_output[3528] = '{87.8344434899};
############ END DEBUG ############*/
test_input[28232:28239] = '{32'hc26074c3, 32'hc11b73e8, 32'hbf6f1b30, 32'h429f24b8, 32'h4084d156, 32'h423a11bc, 32'hc24c70be, 32'h423dc76d};
test_label[3529] = '{32'h423dc76d};
test_output[3529] = '{32'h42008204};
/*############ DEBUG ############
test_input[28232:28239] = '{-56.1140239044, -9.71579780695, -0.934008608224, 79.571718507, 4.15055355186, 46.5173198154, -51.1100992282, 47.4447504908};
test_label[3529] = '{47.4447504908};
test_output[3529] = '{32.1269680163};
############ END DEBUG ############*/
test_input[28240:28247] = '{32'hc296c52c, 32'hc28fae44, 32'hc27075a5, 32'hc0b32e7a, 32'hc2835626, 32'h408e9e7b, 32'hbfc61e43, 32'h421f4da4};
test_label[3530] = '{32'hc2835626};
test_output[3530] = '{32'h42d2fcf8};
/*############ DEBUG ############
test_input[28240:28247] = '{-75.3851049129, -71.8403653622, -60.1148865791, -5.5994236244, -65.6682594369, 4.45684579186, -1.54779845749, 39.8258201075};
test_label[3530] = '{-65.6682594369};
test_output[3530] = '{105.494079544};
############ END DEBUG ############*/
test_input[28248:28255] = '{32'h412439b8, 32'h4285d242, 32'hbfda0494, 32'h414b9936, 32'hc24a2240, 32'hc13ff463, 32'hc2a16b53, 32'hc2c37377};
test_label[3531] = '{32'hc13ff463};
test_output[3531] = '{32'h429dd0ce};
/*############ DEBUG ############
test_input[28248:28255] = '{10.2640915358, 66.910656738, -1.70326470213, 12.7249053039, -50.5334456147, -11.9971643912, -80.7096165547, -97.725513679};
test_label[3531] = '{-11.9971643912};
test_output[3531] = '{78.9078211292};
############ END DEBUG ############*/
test_input[28256:28263] = '{32'hc200bae1, 32'h407d88ab, 32'hc23d9ae9, 32'hc2a2b09a, 32'hc232982b, 32'h42770c32, 32'h428a739a, 32'h40112f03};
test_label[3532] = '{32'h42770c32};
test_output[3532] = '{32'h40eedcc3};
/*############ DEBUG ############
test_input[28256:28263] = '{-32.182499743, 3.96146644106, -47.4012783497, -81.3449243735, -44.6485998069, 61.7619094488, 69.2257848686, 2.26849428693};
test_label[3532] = '{61.7619094488};
test_output[3532] = '{7.4644486851};
############ END DEBUG ############*/
test_input[28264:28271] = '{32'hc27e2f9e, 32'hc2bd5d34, 32'hc2272260, 32'hc1714478, 32'h4290ea1b, 32'hc2410732, 32'h42bfbddf, 32'h42b10e29};
test_label[3533] = '{32'h42b10e29};
test_output[3533] = '{32'h40eb009d};
/*############ DEBUG ############
test_input[28264:28271] = '{-63.5464998083, -94.6820411245, -41.7835676001, -15.0792162858, 72.4572346792, -48.2570256898, 95.8708383135, 88.527660292};
test_label[3533] = '{88.527660292};
test_output[3533] = '{7.34382480345};
############ END DEBUG ############*/
test_input[28272:28279] = '{32'hc2a0baa8, 32'h421d5e12, 32'hc123e905, 32'h4095c4f4, 32'h42c184e9, 32'hc1fc27d4, 32'h41a07d4e, 32'h42aec460};
test_label[3534] = '{32'hc1fc27d4};
test_output[3534] = '{32'h43004774};
/*############ DEBUG ############
test_input[28272:28279] = '{-80.3645599376, 39.3418646136, -10.2443895659, 4.6802922398, 96.7595870579, -31.5194472035, 20.0611839215, 87.3835468972};
test_label[3534] = '{-31.5194472035};
test_output[3534] = '{128.279118988};
############ END DEBUG ############*/
test_input[28280:28287] = '{32'hc19edf54, 32'hc24efb5a, 32'h4298e1d8, 32'hc2c2a758, 32'hc09d8322, 32'h425f7b9e, 32'hc2bf980c, 32'hc1a287cb};
test_label[3535] = '{32'h425f7b9e};
test_output[3535] = '{32'h41a49025};
/*############ DEBUG ############
test_input[28280:28287] = '{-19.8590464237, -51.7454620853, 76.4411015024, -97.3268415163, -4.92225753236, 55.8707189847, -95.7969662495, -20.3163051278};
test_label[3535] = '{55.8707189847};
test_output[3535] = '{20.5703825189};
############ END DEBUG ############*/
test_input[28288:28295] = '{32'hc09dcb1d, 32'h42b2675b, 32'hc1b7c632, 32'h429299d5, 32'hc2a77c98, 32'hc286fe25, 32'h4232dc14, 32'hc2b26230};
test_label[3536] = '{32'hc1b7c632};
test_output[3536] = '{32'h42e058e7};
/*############ DEBUG ############
test_input[28288:28295] = '{-4.9310442061, 89.2018639902, -22.9717749167, 73.3004522124, -83.7433481582, -67.4963785596, 44.7149198534, -89.1917756138};
test_label[3536] = '{-22.9717749167};
test_output[3536] = '{112.173639031};
############ END DEBUG ############*/
test_input[28296:28303] = '{32'h42aeae80, 32'hc0a74b7d, 32'h42314195, 32'hbfd72f39, 32'hc18a3ab6, 32'hc2a54fd8, 32'h426e2989, 32'hc2a54e9a};
test_label[3537] = '{32'hc2a54e9a};
test_output[3537] = '{32'h4329fe8d};
/*############ DEBUG ############
test_input[28296:28303] = '{87.3408168847, -5.22796466373, 44.3140431392, -1.6811286694, -17.2786670473, -82.6559437516, 59.5405599749, -82.6535189686};
test_label[3537] = '{-82.6535189686};
test_output[3537] = '{169.994335853};
############ END DEBUG ############*/
test_input[28304:28311] = '{32'hc2b65444, 32'h420d58e5, 32'h41dbbb77, 32'hc191ec3f, 32'hc2c05d59, 32'h41864091, 32'h41c7d229, 32'h424f7aeb};
test_label[3538] = '{32'h424f7aeb};
test_output[3538] = '{32'h338dd8ed};
/*############ DEBUG ############
test_input[28304:28311] = '{-91.1645803076, 35.3368123575, 27.4665364699, -18.2403551383, -96.1823177738, 16.7815257893, 24.9776172096, 51.8700368415};
test_label[3538] = '{51.8700368415};
test_output[3538] = '{6.60528297224e-08};
############ END DEBUG ############*/
test_input[28312:28319] = '{32'h42098a21, 32'hc28b557d, 32'h419bb113, 32'hc1718ff7, 32'h42739277, 32'hc219086a, 32'h425c9a58, 32'hc2847970};
test_label[3539] = '{32'hc1718ff7};
test_output[3539] = '{32'h4297fcde};
/*############ DEBUG ############
test_input[28312:28319] = '{34.3848908595, -69.666968309, 19.4614619604, -15.0976477225, 60.8930326696, -38.258217953, 55.1507252093, -66.2371854238};
test_label[3539] = '{-15.0976477225};
test_output[3539] = '{75.9938826184};
############ END DEBUG ############*/
test_input[28320:28327] = '{32'h41a77c14, 32'h423b96b7, 32'h424252e2, 32'hc243b002, 32'h410c45d3, 32'h426dff6c, 32'hc1ff841e, 32'h427b6382};
test_label[3540] = '{32'h424252e2};
test_output[3540] = '{32'h4164d00f};
/*############ DEBUG ############
test_input[28320:28327] = '{20.9355849305, 46.8971818027, 48.5809394894, -48.9218812954, 8.76704675937, 59.4994349148, -31.9395110779, 62.8471745896};
test_label[3540] = '{48.5809394894};
test_output[3540] = '{14.3007954528};
############ END DEBUG ############*/
test_input[28328:28335] = '{32'hc281e20b, 32'hc23ab8b9, 32'h42ab9636, 32'hc1b311a8, 32'hc2bd280f, 32'h42b66ef8, 32'hc19b9c7e, 32'h42bef835};
test_label[3541] = '{32'hc281e20b};
test_output[3541] = '{32'h432070b4};
/*############ DEBUG ############
test_input[28328:28335] = '{-64.9414865048, -46.6803947487, 85.7933836082, -22.3836221077, -94.5782398639, 91.2167344293, -19.4514113607, 95.4847805913};
test_label[3541] = '{-64.9414865048};
test_output[3541] = '{160.44023996};
############ END DEBUG ############*/
test_input[28336:28343] = '{32'h42b11da1, 32'h41cfcba4, 32'h426052b6, 32'hc1add193, 32'hc2b58a41, 32'hc27e39da, 32'hc1de9ebc, 32'h424afa2a};
test_label[3542] = '{32'hc1add193};
test_output[3542] = '{32'h42dc9205};
/*############ DEBUG ############
test_input[28336:28343] = '{88.5578656254, 25.9744344898, 56.0807726743, -21.72733047, -90.7700308131, -63.5564951654, -27.8275063595, 50.7443011121};
test_label[3542] = '{-21.72733047};
test_output[3542] = '{110.285196095};
############ END DEBUG ############*/
test_input[28344:28351] = '{32'h4155f885, 32'hc1ec73ee, 32'h429b8350, 32'h41fdf54b, 32'h4282cc13, 32'hc286b95f, 32'hc289401d, 32'hc29da831};
test_label[3543] = '{32'h41fdf54b};
test_output[3543] = '{32'h42380bfb};
/*############ DEBUG ############
test_input[28344:28351] = '{13.3731736979, -29.5566069419, 77.7564677858, 31.7447725855, 65.3985811593, -67.3620527162, -68.6252201994, -78.8285017204};
test_label[3543] = '{31.7447725855};
test_output[3543] = '{46.0116994961};
############ END DEBUG ############*/
test_input[28352:28359] = '{32'hc11d2cde, 32'hc2708cb5, 32'h42bc9e9b, 32'h420f50ec, 32'hc28dea80, 32'hc249049d, 32'h429d9bed, 32'h425a93c1};
test_label[3544] = '{32'hc249049d};
test_output[3544] = '{32'h43109075};
/*############ DEBUG ############
test_input[28352:28359] = '{-9.82345419798, -60.1374098156, 94.3097793323, 35.8290259223, -70.9580043116, -50.2545056458, 78.8045411426, 54.6442925495};
test_label[3544] = '{-50.2545056458};
test_output[3544] = '{144.564285163};
############ END DEBUG ############*/
test_input[28360:28367] = '{32'h422565ee, 32'hc2a6d8f9, 32'h4271d50a, 32'h421831d8, 32'h41cca1a4, 32'hbf8610cd, 32'hc182b035, 32'hc22f99cd};
test_label[3545] = '{32'hc2a6d8f9};
test_output[3545] = '{32'h430fe1bf};
/*############ DEBUG ############
test_input[28360:28367] = '{41.3495402307, -83.4237736114, 60.4580458863, 38.0486769721, 25.5789255616, -1.04738766489, -16.3360393832, -43.9001954315};
test_label[3545] = '{-83.4237736114};
test_output[3545] = '{143.881819503};
############ END DEBUG ############*/
test_input[28368:28375] = '{32'h42ba4ed4, 32'h429b275b, 32'h4120c07f, 32'hc2bfebbf, 32'hc2343f7f, 32'hc2b42f12, 32'h426c1bf4, 32'h418f5fb8};
test_label[3546] = '{32'h426c1bf4};
test_output[3546] = '{32'h420881b3};
/*############ DEBUG ############
test_input[28368:28375] = '{93.1539579845, 77.5768654339, 10.0469963032, -95.9604449267, -45.0620097023, -90.091932129, 59.0272977501, 17.9217376415};
test_label[3546] = '{59.0272977501};
test_output[3546] = '{34.1266604061};
############ END DEBUG ############*/
test_input[28376:28383] = '{32'hc286b739, 32'h42b2a86f, 32'hc28c0160, 32'hc15fff2c, 32'hc285d030, 32'h4242fc58, 32'hc169b627, 32'hc19d1c29};
test_label[3547] = '{32'hc286b739};
test_output[3547] = '{32'h431cafd4};
/*############ DEBUG ############
test_input[28376:28383] = '{-67.3578587509, 89.3289695456, -70.0026854296, -13.9997981461, -66.9066148811, 48.7464307863, -14.6069710305, -19.6387508685};
test_label[3547] = '{-67.3578587509};
test_output[3547] = '{156.686828297};
############ END DEBUG ############*/
test_input[28384:28391] = '{32'hc2a19a34, 32'hc1ec92a5, 32'h4298e2b4, 32'hc172de09, 32'h4275243c, 32'h402d3e53, 32'hc0c8a72e, 32'h42a55549};
test_label[3548] = '{32'h402d3e53};
test_output[3548] = '{32'h429fec5a};
/*############ DEBUG ############
test_input[28384:28391] = '{-80.8011809128, -29.5716042132, 76.4427804025, -15.1792080759, 61.2853839539, 2.70692887478, -6.27040787355, 82.6665731672};
test_label[3548] = '{2.70692887478};
test_output[3548] = '{79.9616240467};
############ END DEBUG ############*/
test_input[28392:28399] = '{32'hc2731aaa, 32'hc26953b5, 32'hc150b242, 32'h41c6148e, 32'h429d7883, 32'h4288a649, 32'hc19f91e0, 32'h42ba0e2b};
test_label[3549] = '{32'h42ba0e2b};
test_output[3549] = '{32'h3526a4ab};
/*############ DEBUG ############
test_input[28392:28399] = '{-60.7760379847, -58.3317460718, -13.043520268, 24.7600367512, 78.7353744311, 68.3247720389, -19.946228972, 93.0276701056};
test_label[3549] = '{93.0276701056};
test_output[3549] = '{6.20794409281e-07};
############ END DEBUG ############*/
test_input[28400:28407] = '{32'hc212ee10, 32'hc2c54f5f, 32'h42146298, 32'hc280ef9e, 32'hc01cce72, 32'hc20f1131, 32'hc295bf3e, 32'h4227e0fa};
test_label[3550] = '{32'hc212ee10};
test_output[3550] = '{32'h429d6b6b};
/*############ DEBUG ############
test_input[28400:28407] = '{-36.7324837844, -98.6550244024, 37.0962817033, -64.467998645, -2.45010042231, -35.7667899927, -74.8735185721, 41.9697020116};
test_label[3550] = '{-36.7324837844};
test_output[3550] = '{78.7098038696};
############ END DEBUG ############*/
test_input[28408:28415] = '{32'h413f42ba, 32'h40ac055f, 32'hc2a98669, 32'hc2a7dc13, 32'hc297d695, 32'h425fad0c, 32'hc283183e, 32'h423a6bbb};
test_label[3551] = '{32'hc2a98669};
test_output[3551] = '{32'h430cae7d};
/*############ DEBUG ############
test_input[28408:28415] = '{11.9537908916, 5.37565557543, -84.7625194655, -83.9298340192, -75.9191037079, 55.9189911571, -65.5473512088, 46.6052046221};
test_label[3551] = '{-84.7625194655};
test_output[3551] = '{140.681600791};
############ END DEBUG ############*/
test_input[28416:28423] = '{32'h4281f56b, 32'hc2818180, 32'hc2b656a1, 32'hc25539c8, 32'hc2b386d0, 32'hc1f1914f, 32'h40301faa, 32'h41f46e5b};
test_label[3552] = '{32'h41f46e5b};
test_output[3552] = '{32'h4209b3a8};
/*############ DEBUG ############
test_input[28416:28423] = '{64.9793294061, -64.7529313661, -91.169199766, -53.3064276763, -89.7633065234, -30.1959506062, 2.75193270481, 30.5538838263};
test_label[3552] = '{30.5538838263};
test_output[3552] = '{34.4254455798};
############ END DEBUG ############*/
test_input[28424:28431] = '{32'hc1440386, 32'hc0a49714, 32'h41fb448f, 32'hc2bb767b, 32'hc08e6b59, 32'h4220db07, 32'hc2a52be4, 32'hc29dae1a};
test_label[3553] = '{32'h41fb448f};
test_output[3553] = '{32'h410ce399};
/*############ DEBUG ############
test_input[28424:28431] = '{-12.2508605201, -5.1434422275, 31.4084764413, -93.7314058433, -4.45060382829, 40.2138928064, -82.5857254167, -78.8400402576};
test_label[3553] = '{31.4084764413};
test_output[3553] = '{8.80556627271};
############ END DEBUG ############*/
test_input[28432:28439] = '{32'h417f3d2e, 32'h426791eb, 32'h420f07e3, 32'hbf9ca04d, 32'h4286fe0b, 32'hc2bdcc1a, 32'h429291cb, 32'h42ba7671};
test_label[3554] = '{32'hbf9ca04d};
test_output[3554] = '{32'h42bce8f2};
/*############ DEBUG ############
test_input[28432:28439] = '{15.9524363014, 57.8924991644, 35.7577015741, -1.2236419427, 67.4961742884, -94.898634471, 73.284754532, 93.2313270831};
test_label[3554] = '{-1.2236419427};
test_output[3554] = '{94.454969028};
############ END DEBUG ############*/
test_input[28440:28447] = '{32'h40761a0c, 32'h423fbd89, 32'hc16479d0, 32'h42b80d64, 32'h4253a8ae, 32'hc1f2f7fe, 32'h42a4bf18, 32'hc2471c42};
test_label[3555] = '{32'h40761a0c};
test_output[3555] = '{32'h42b05c9c};
/*############ DEBUG ############
test_input[28440:28447] = '{3.84533971276, 47.9350912885, -14.2797396101, 92.0261500462, 52.9147280118, -30.3710900437, 82.3732278692, -49.7775946764};
test_label[3555] = '{3.84533971276};
test_output[3555] = '{88.1808745689};
############ END DEBUG ############*/
test_input[28448:28455] = '{32'hc0f898e7, 32'h42b87437, 32'h42a05a67, 32'h41c7bcf9, 32'h424df289, 32'h4276d8f8, 32'h40bda545, 32'hc28a8e7f};
test_label[3556] = '{32'hc28a8e7f};
test_output[3556] = '{32'h4321815b};
/*############ DEBUG ############
test_input[28448:28455] = '{-7.76866494507, 92.2269792148, 80.1765660634, 24.9672716652, 51.4868520241, 61.7118817756, 5.92642427473, -69.2783100871};
test_label[3556] = '{-69.2783100871};
test_output[3556] = '{161.505295144};
############ END DEBUG ############*/
test_input[28456:28463] = '{32'hc2b6c4d3, 32'hc291ec12, 32'h41cf2737, 32'hc298aa9c, 32'h41dae565, 32'h42a59ee8, 32'hc28c43d6, 32'h426e874f};
test_label[3557] = '{32'hc291ec12};
test_output[3557] = '{32'h431bc57d};
/*############ DEBUG ############
test_input[28456:28463] = '{-91.3844241595, -72.9610763986, 25.8941487966, -76.3332240744, 27.3620097816, 82.8103662501, -70.1324947894, 59.6321373288};
test_label[3557] = '{-72.9610763986};
test_output[3557] = '{155.771442649};
############ END DEBUG ############*/
test_input[28464:28471] = '{32'hc2abf8cb, 32'hc031d795, 32'h41b0c12e, 32'hc2837404, 32'h411b0573, 32'hc28cca35, 32'hc2311691, 32'hc2368dc4};
test_label[3558] = '{32'hc2837404};
test_output[3558] = '{32'h42afa450};
/*############ DEBUG ############
test_input[28464:28471] = '{-85.985920614, -2.77878308219, 22.0943264077, -65.7265944535, 9.68882991633, -70.3949390751, -44.272038665, -45.6384437944};
test_label[3558] = '{-65.7265944535};
test_output[3558] = '{87.8209249573};
############ END DEBUG ############*/
test_input[28472:28479] = '{32'hc26cf9c8, 32'h4228498e, 32'h42b417d4, 32'h4296bc44, 32'hc2c490af, 32'hc2515e2c, 32'h4207c951, 32'h41f074bb};
test_label[3559] = '{32'h4207c951};
test_output[3559] = '{32'h42606658};
/*############ DEBUG ############
test_input[28472:28479] = '{-59.2439285647, 42.0718314802, 90.0465420438, 75.3677070575, -98.2825877807, -52.3419664197, 33.9465990676, 30.0569965975};
test_label[3559] = '{33.9465990676};
test_output[3559] = '{56.099943398};
############ END DEBUG ############*/
test_input[28480:28487] = '{32'hc1f1d91c, 32'h429e7da1, 32'h41f9eca3, 32'hc18e1d94, 32'h428c9cf1, 32'h4287e1f4, 32'h41eddd0f, 32'h4207ec8e};
test_label[3560] = '{32'h4207ec8e};
test_output[3560] = '{32'h42350eda};
/*############ DEBUG ############
test_input[28480:28487] = '{-30.2310105887, 79.2453693203, 31.2405461984, -17.7644430762, 70.3065238872, 67.9413128362, 29.7329391175, 33.9810095036};
test_label[3560] = '{33.9810095036};
test_output[3560] = '{45.2645033216};
############ END DEBUG ############*/
test_input[28488:28495] = '{32'h42bc927f, 32'hc29f61a9, 32'h41ecce1f, 32'h41ebd7f1, 32'hc204844b, 32'h3ee87f30, 32'hc28cd1bc, 32'hc26778fb};
test_label[3561] = '{32'h41ebd7f1};
test_output[3561] = '{32'h42819c82};
/*############ DEBUG ############
test_input[28488:28495] = '{94.2861233289, -79.6907419295, 29.6006452346, 29.4804408701, -33.1291926816, 0.454095355434, -70.4096346758, -57.868143368};
test_label[3561] = '{29.4804408701};
test_output[3561] = '{64.8056824588};
############ END DEBUG ############*/
test_input[28496:28503] = '{32'h42573bd3, 32'h42816bb8, 32'h42593d3c, 32'h4268c97a, 32'hc15a88b3, 32'h418bf129, 32'hc20c99a8, 32'hc2ac2808};
test_label[3562] = '{32'hc20c99a8};
test_output[3562] = '{32'h42c7b955};
/*############ DEBUG ############
test_input[28496:28503] = '{53.8084224705, 64.7103903477, 54.3097993859, 58.1967540938, -13.6583735025, 17.4927547199, -35.1500531243, -86.0781888701};
test_label[3562] = '{-35.1500531243};
test_output[3562] = '{99.8619742134};
############ END DEBUG ############*/
test_input[28504:28511] = '{32'hc18567d2, 32'h42b9ba34, 32'h41d9e0af, 32'hc1ada872, 32'h4124f196, 32'hc23e25a8, 32'hc0ffd202, 32'h423ab072};
test_label[3563] = '{32'h4124f196};
test_output[3563] = '{32'h42a51c01};
/*############ DEBUG ############
test_input[28504:28511] = '{-16.6756933713, 92.8636795418, 27.2347084862, -21.7072485583, 10.3089809985, -47.5367726832, -7.99438584358, 46.6723112085};
test_label[3563] = '{10.3089809985};
test_output[3563] = '{82.5546985433};
############ END DEBUG ############*/
test_input[28512:28519] = '{32'hc28d1e2f, 32'hc12cf372, 32'h403e0bb3, 32'hc220106d, 32'h42b3267d, 32'h4259bf58, 32'hc0a956e1, 32'h42154974};
test_label[3564] = '{32'hc28d1e2f};
test_output[3564] = '{32'h43202256};
/*############ DEBUG ############
test_input[28512:28519] = '{-70.5589505014, -10.809434696, 2.96946408067, -40.0160425329, 89.5751757835, 54.4368577464, -5.29185556595, 37.3217324498};
test_label[3564] = '{-70.5589505014};
test_output[3564] = '{160.134126285};
############ END DEBUG ############*/
test_input[28520:28527] = '{32'h429048e8, 32'hc1a5940f, 32'hc2215a4f, 32'h41d8ed83, 32'h42428bf4, 32'hc2a29c3e, 32'h4238c65b, 32'h4233e2ee};
test_label[3565] = '{32'h4233e2ee};
test_output[3565] = '{32'h41d95dc5};
/*############ DEBUG ############
test_input[28520:28527] = '{72.1423985293, -20.6972951545, -40.3381932078, 27.1159734376, 48.636673776, -81.3051606948, 46.1937054875, 44.9716128838};
test_label[3565] = '{44.9716128838};
test_output[3565] = '{27.1707856456};
############ END DEBUG ############*/
test_input[28528:28535] = '{32'h429bac7e, 32'h3eb03d35, 32'h42557127, 32'h428390f9, 32'h424ff761, 32'hc2019cc2, 32'h4291dafa, 32'hc0b5d23b};
test_label[3566] = '{32'hc0b5d23b};
test_output[3566] = '{32'h42a70d65};
/*############ DEBUG ############
test_input[28528:28535] = '{77.8368951211, 0.344216986407, 53.3605019074, 65.7831530276, 51.9915814095, -32.403085379, 72.9276900652, -5.6819127375};
test_label[3566] = '{-5.6819127375};
test_output[3566] = '{83.5261649032};
############ END DEBUG ############*/
test_input[28536:28543] = '{32'hc278f748, 32'hc21fd368, 32'hc2b0ffa0, 32'hc29ace03, 32'h4289cda2, 32'hc201c049, 32'h42706dea, 32'hc24cb294};
test_label[3567] = '{32'hc24cb294};
test_output[3567] = '{32'h42f02700};
/*############ DEBUG ############
test_input[28536:28543] = '{-62.2414857915, -39.9564530859, -88.4992709894, -77.4023651818, 68.9016242611, -32.4377770469, 60.1073380534, -51.1743934821};
test_label[3567] = '{-51.1743934821};
test_output[3567] = '{120.076169329};
############ END DEBUG ############*/
test_input[28544:28551] = '{32'hc293ccf2, 32'hc2a751c1, 32'h426599d6, 32'h41ba8f77, 32'hc1d305d6, 32'hc27ea04d, 32'hc2455462, 32'h429a7d33};
test_label[3568] = '{32'h41ba8f77};
test_output[3568] = '{32'h4257b2aa};
/*############ DEBUG ############
test_input[28544:28551] = '{-73.9002848359, -83.6596749654, 57.4002300073, 23.3200519746, -26.3778492484, -63.6565434433, -49.332405623, 77.2445274095};
test_label[3568] = '{23.3200519746};
test_output[3568] = '{53.9244754373};
############ END DEBUG ############*/
test_input[28552:28559] = '{32'h41a759a4, 32'h4265ce99, 32'h4083670d, 32'hc23d8ce1, 32'h42ba1082, 32'hc1c51d7c, 32'h422c2d88, 32'h424c753c};
test_label[3569] = '{32'h422c2d88};
test_output[3569] = '{32'h4247f37b};
/*############ DEBUG ############
test_input[28552:28559] = '{20.9187695882, 57.4517541631, 4.10632938408, -47.3875774842, 93.032238271, -24.6393970141, 43.0444651529, 51.1144875247};
test_label[3569] = '{43.0444651529};
test_output[3569] = '{49.9877731181};
############ END DEBUG ############*/
test_input[28560:28567] = '{32'hc1f184c9, 32'h423c496c, 32'h42172284, 32'hc2ab9429, 32'hc2b65ec0, 32'hc28b91bd, 32'hbf678fb5, 32'hc255c490};
test_label[3570] = '{32'hc1f184c9};
test_output[3570] = '{32'h429a85f4};
/*############ DEBUG ############
test_input[28560:28567] = '{-30.1898364253, 47.0717001854, 37.7837077445, -85.789378295, -91.1850580698, -69.7846477035, -0.904536565578, -53.4419538796};
test_label[3570] = '{-30.1898364253};
test_output[3570] = '{77.2616291351};
############ END DEBUG ############*/
test_input[28568:28575] = '{32'hc2c653cc, 32'hc229172f, 32'h4146c76e, 32'hc17cbb37, 32'h41e11b0d, 32'hc25fb231, 32'h4218682f, 32'hc2a923ad};
test_label[3571] = '{32'h4218682f};
test_output[3571] = '{32'h38457d05};
/*############ DEBUG ############
test_input[28568:28575] = '{-99.1636628083, -42.2726396508, 12.4236885323, -15.7957070425, 28.1382082204, -55.92401396, 38.1017431849, -84.5696787064};
test_label[3571] = '{38.1017431849};
test_output[3571] = '{4.70848927258e-05};
############ END DEBUG ############*/
test_input[28576:28583] = '{32'h41c12afd, 32'h428e3c97, 32'h42bfa884, 32'h41d5224a, 32'h42b39a61, 32'h42a4d5d4, 32'hc26eb1a6, 32'h42255416};
test_label[3572] = '{32'h42bfa884};
test_output[3572] = '{32'h3b1dee5d};
/*############ DEBUG ############
test_input[28576:28583] = '{24.1459894272, 71.1183409477, 95.8291353245, 26.6417433886, 89.8015235163, 82.4176317596, -59.6734862626, 41.3321140473};
test_label[3572] = '{95.8291353245};
test_output[3572] = '{0.00240983746568};
############ END DEBUG ############*/
test_input[28584:28591] = '{32'hc28c1ca1, 32'hc24bdf66, 32'h4294b31f, 32'h42917c74, 32'hc2970f82, 32'hc27f2920, 32'h4294f2a8, 32'h4223dd00};
test_label[3573] = '{32'h4294b31f};
test_output[3573] = '{32'h3f58d52d};
/*############ DEBUG ############
test_input[28584:28591] = '{-70.0559132898, -50.9681610416, 74.3498491257, 72.7430706246, -75.5302898228, -63.7901607402, 74.4739344156, 40.9658199777};
test_label[3573] = '{74.3498491257};
test_output[3573] = '{0.847002823153};
############ END DEBUG ############*/
test_input[28592:28599] = '{32'h41e6cfdb, 32'hc2306266, 32'hc253cd0f, 32'hc1a198dc, 32'h42a6eace, 32'h42b3c34d, 32'hc290335a, 32'hc1d6c928};
test_label[3574] = '{32'hc1d6c928};
test_output[3574] = '{32'h42e9766b};
/*############ DEBUG ############
test_input[28592:28599] = '{28.8514928546, -44.0960918286, -52.9502538886, -20.199638734, 83.4586046618, 89.8814437247, -72.1002922414, -26.8482210761};
test_label[3574] = '{-26.8482210761};
test_output[3574] = '{116.731287522};
############ END DEBUG ############*/
test_input[28600:28607] = '{32'h42b545b6, 32'hc1f69238, 32'hc2b0b621, 32'hc20cd7c5, 32'h4211ba66, 32'hc259e463, 32'h40ab091d, 32'hc2c03fb9};
test_label[3575] = '{32'h4211ba66};
test_output[3575] = '{32'h4258d106};
/*############ DEBUG ############
test_input[28600:28607] = '{90.6361560705, -30.8213967279, -88.3557201762, -35.2107140697, 36.4320301519, -54.4730337995, 5.34486265974, -96.1244574481};
test_label[3575] = '{36.4320301519};
test_output[3575] = '{54.2041259186};
############ END DEBUG ############*/
test_input[28608:28615] = '{32'h414525db, 32'h42ac8206, 32'hc2148213, 32'h419a25c2, 32'h4198bbc7, 32'h40af58b4, 32'hc2711a6e, 32'hc0d23509};
test_label[3576] = '{32'hc2711a6e};
test_output[3576] = '{32'h4312879e};
/*############ DEBUG ############
test_input[28608:28615] = '{12.3217422236, 86.2539529744, -37.1270244429, 19.2684370589, 19.0916874596, 5.47957784654, -60.275808887, -6.56897383745};
test_label[3576] = '{-60.275808887};
test_output[3576] = '{146.529761861};
############ END DEBUG ############*/
test_input[28616:28623] = '{32'h42a4db43, 32'hc1a05b58, 32'h4272c02f, 32'h4253a91b, 32'h40f28afe, 32'h4284a72f, 32'hc173e32e, 32'hc1274a42};
test_label[3577] = '{32'h42a4db43};
test_output[3577] = '{32'h33db1278};
/*############ DEBUG ############
test_input[28616:28623] = '{82.4282454542, -20.0446016941, 60.6876803284, 52.9151410099, 7.57946703356, 66.3265318436, -15.2429637226, -10.455629385};
test_label[3577] = '{82.4282454542};
test_output[3577] = '{1.02013413369e-07};
############ END DEBUG ############*/
test_input[28624:28631] = '{32'hc22ee420, 32'hc23c8d1b, 32'h42c23be7, 32'hc2b5bb07, 32'h429ec7cc, 32'hc28110cb, 32'hc2c28a1c, 32'hc1c604ab};
test_label[3578] = '{32'hc1c604ab};
test_output[3578] = '{32'h42f3bd11};
/*############ DEBUG ############
test_input[28624:28631] = '{-43.7227778114, -47.1377985006, 97.1169931361, -90.8652856884, 79.390227773, -64.5328006228, -97.2697437796, -24.7522786722};
test_label[3578] = '{-24.7522786722};
test_output[3578] = '{121.869271828};
############ END DEBUG ############*/
test_input[28632:28639] = '{32'h4189ece0, 32'hc287337d, 32'h420b0378, 32'hc18d2998, 32'h410d67f4, 32'hc21c1504, 32'hc25b9281, 32'h424f149a};
test_label[3579] = '{32'hc287337d};
test_output[3579] = '{32'h42eebdca};
/*############ DEBUG ############
test_input[28632:28639] = '{17.240661704, -67.6005661861, 34.7533885797, -17.6453086523, 8.83787939598, -39.0205246204, -54.8930688732, 51.7701168688};
test_label[3579] = '{-67.6005661861};
test_output[3579] = '{119.370683096};
############ END DEBUG ############*/
test_input[28640:28647] = '{32'h423c0069, 32'h4295068c, 32'hc29fba14, 32'hc2a55d40, 32'hc2bdb3d8, 32'h425083c6, 32'hc25ccdf1, 32'hc268eb55};
test_label[3580] = '{32'h425083c6};
test_output[3580] = '{32'h41b312a5};
/*############ DEBUG ############
test_input[28640:28647] = '{47.0003988397, 74.5127902712, -79.8634368004, -82.6821293557, -94.8512541978, 52.1286867987, -55.2011147213, -58.2298164045};
test_label[3580] = '{52.1286867987};
test_output[3580] = '{22.3841034726};
############ END DEBUG ############*/
test_input[28648:28655] = '{32'h4082ca0f, 32'h424cd9ea, 32'h4175707f, 32'hc289938c, 32'hc0a3508e, 32'hc2b745a8, 32'hc2c17361, 32'h42a6c164};
test_label[3581] = '{32'hc0a3508e};
test_output[3581] = '{32'h42b0f66d};
/*############ DEBUG ############
test_input[28648:28655] = '{4.08716555748, 51.212804952, 15.3399653262, -68.7881799505, -5.1035832964, -91.6360502507, -96.7253521841, 83.3777166673};
test_label[3581] = '{-5.1035832964};
test_output[3581] = '{88.4812999637};
############ END DEBUG ############*/
test_input[28656:28663] = '{32'hc1f07fd5, 32'h427dae82, 32'h429df7aa, 32'hc254336f, 32'hc25362dc, 32'h424a2b8f, 32'hc214c8d3, 32'h429054a7};
test_label[3582] = '{32'h429df7aa};
test_output[3582] = '{32'h3a8f4548};
/*############ DEBUG ############
test_input[28656:28663] = '{-30.062418342, 63.4204166587, 78.9837178015, -53.0502282985, -52.8465428293, 50.54253721, -37.1961155447, 72.1653384496};
test_label[3582] = '{78.9837178015};
test_output[3582] = '{0.00109306819412};
############ END DEBUG ############*/
test_input[28664:28671] = '{32'h424adf87, 32'h40302c08, 32'h429a7c4b, 32'h42c251bc, 32'hc27a2cd4, 32'h42c4521d, 32'hc1cfff94, 32'hc0edd8d0};
test_label[3583] = '{32'h42c4521d};
test_output[3583] = '{32'h3ea049c7};
/*############ DEBUG ############
test_input[28664:28671] = '{50.7182901119, 2.75268735644, 77.2427601425, 97.1596371, -62.5437773702, 98.1603765898, -25.999793844, -7.43271643264};
test_label[3583] = '{98.1603765898};
test_output[3583] = '{0.313062862432};
############ END DEBUG ############*/
test_input[28672:28679] = '{32'hc27a3712, 32'h418b7926, 32'hc0a8cf60, 32'h42326c18, 32'h426c3e6b, 32'hc12b8c42, 32'hc1dfaed0, 32'hc1a24cb9};
test_label[3584] = '{32'hc27a3712};
test_output[3584] = '{32'h42f33abe};
/*############ DEBUG ############
test_input[28672:28679] = '{-62.5537792908, 17.434155413, -5.27531414505, 44.6055602298, 59.0609538744, -10.7217426918, -27.9603571822, -20.2874620361};
test_label[3584] = '{-62.5537792908};
test_output[3584] = '{121.614733693};
############ END DEBUG ############*/
test_input[28680:28687] = '{32'h42a22d29, 32'h424e3bab, 32'h41f23d38, 32'h4289bc98, 32'h42804b8d, 32'hc09b7e34, 32'h427aa9dd, 32'hc28dd7a1};
test_label[3585] = '{32'hc09b7e34};
test_output[3585] = '{32'h42abe50d};
/*############ DEBUG ############
test_input[28680:28687] = '{81.0882010824, 51.5582711408, 30.2798920234, 68.868343748, 64.1475595373, -4.85915579991, 62.6658809825, -70.9211513957};
test_label[3585] = '{-4.85915579991};
test_output[3585] = '{85.9473618677};
############ END DEBUG ############*/
test_input[28688:28695] = '{32'hc22dcda7, 32'hc22e1e74, 32'h41ea51e0, 32'hc15a81aa, 32'h413fd7ea, 32'hc2c7db04, 32'hc275acae, 32'h41a2e8fb};
test_label[3586] = '{32'h413fd7ea};
test_output[3586] = '{32'h418a6630};
/*############ DEBUG ############
test_input[28688:28695] = '{-43.4508324171, -43.5297374988, 29.289977437, -13.656655821, 11.9902137103, -99.9277621535, -61.4186342735, 20.3637599187};
test_label[3586] = '{11.9902137103};
test_output[3586] = '{17.2998966082};
############ END DEBUG ############*/
test_input[28696:28703] = '{32'h41c44f1a, 32'hc272d445, 32'h42b5cb9f, 32'hc27d402c, 32'hc2b7f2ba, 32'hc28b9d6f, 32'hc2b1f15b, 32'hc2c7f384};
test_label[3587] = '{32'h42b5cb9f};
test_output[3587] = '{32'h80000000};
/*############ DEBUG ############
test_input[28696:28703] = '{24.5386235027, -60.7072938485, 90.8976973797, -63.3126688178, -91.9740727913, -69.8074859951, -88.9713966217, -99.9756161403};
test_label[3587] = '{90.8976973797};
test_output[3587] = '{-0.0};
############ END DEBUG ############*/
test_input[28704:28711] = '{32'hc26360ea, 32'h42a5e8ea, 32'h41cebe94, 32'hc20cfad6, 32'hc280b323, 32'h40d2aa4a, 32'hc1fc1fa4, 32'hc197414f};
test_label[3588] = '{32'h41cebe94};
test_output[3588] = '{32'h42647289};
/*############ DEBUG ############
test_input[28704:28711] = '{-56.8446429154, 82.9549073329, 25.8430554561, -35.2449566972, -64.3498794358, 6.5832870713, -31.5154502722, -18.9068884324};
test_label[3588] = '{25.8430554561};
test_output[3588] = '{57.1118518768};
############ END DEBUG ############*/
test_input[28712:28719] = '{32'hc2835e36, 32'hc19c111a, 32'hc250ae2f, 32'h418c4b2b, 32'h41c68624, 32'hc1e93276, 32'hc2b3e05a, 32'h423b5e18};
test_label[3589] = '{32'hc2b3e05a};
test_output[3589] = '{32'h4308c7b3};
/*############ DEBUG ############
test_input[28712:28719] = '{-65.6840080788, -19.5083507531, -52.1701016935, 17.5367032409, 24.8154988167, -29.1496397592, -89.9381842006, 46.8418871203};
test_label[3589] = '{-89.9381842006};
test_output[3589] = '{136.780071321};
############ END DEBUG ############*/
test_input[28720:28727] = '{32'h410f3c98, 32'h41e289d7, 32'hc1090191, 32'hc2166779, 32'hc029550b, 32'h42b72f8f, 32'h42a8dd96, 32'h42bfa7dd};
test_label[3590] = '{32'h410f3c98};
test_output[3590] = '{32'h42adc7a7};
/*############ DEBUG ############
test_input[28720:28727] = '{8.95229348822, 28.3173053015, -8.56288257365, -37.6010482207, -2.64581554056, 91.5928854279, 84.4327888207, 95.8278556185};
test_label[3590] = '{8.95229348822};
test_output[3590] = '{86.8899496248};
############ END DEBUG ############*/
test_input[28728:28735] = '{32'hc2c1aa25, 32'h419451e9, 32'h41975010, 32'h42ae19e0, 32'hc2b708de, 32'hc26e349d, 32'hc2c15605, 32'h42b7c589};
test_label[3591] = '{32'h42ae19e0};
test_output[3591] = '{32'h409afb64};
/*############ DEBUG ############
test_input[28728:28735] = '{-96.8323098998, 18.5399949907, 18.9140939338, 87.0505395521, -91.5173187475, -59.5513784501, -96.6680040839, 91.8858139243};
test_label[3591] = '{87.0505395521};
test_output[3591] = '{4.84318748904};
############ END DEBUG ############*/
test_input[28736:28743] = '{32'h42c4dc3a, 32'h4250fee8, 32'h41fa98cb, 32'h42a6538a, 32'hc2a38b38, 32'h42903769, 32'h42a94832, 32'h42b3abe0};
test_label[3592] = '{32'h4250fee8};
test_output[3592] = '{32'h4238b9be};
/*############ DEBUG ############
test_input[28736:28743] = '{98.4301320678, 52.2489313415, 31.3246059587, 83.1631659696, -81.7719142479, 72.1082243717, 84.6410089092, 89.8356956753};
test_label[3592] = '{52.2489313415};
test_output[3592] = '{46.1813871029};
############ END DEBUG ############*/
test_input[28744:28751] = '{32'hc1ad77a6, 32'h4212ac06, 32'hc15c007e, 32'hc0c04215, 32'h425407bb, 32'hc283622f, 32'h425e3261, 32'hc0f2f715};
test_label[3593] = '{32'hc283622f};
test_output[3593] = '{32'h42f2a22d};
/*############ DEBUG ############
test_input[28744:28751] = '{-21.6834218917, 36.6679905324, -13.7501204915, -6.00806682451, 53.0075484908, -65.6917639421, 55.5491982668, -7.59266158618};
test_label[3593] = '{-65.6917639421};
test_output[3593] = '{121.316752566};
############ END DEBUG ############*/
test_input[28752:28759] = '{32'hc0ae2ad8, 32'h41913b3c, 32'h41b63fe5, 32'hc2bdba3c, 32'hc22cec5f, 32'h42c7b1f3, 32'h42917ad3, 32'h42ab605e};
test_label[3594] = '{32'hc22cec5f};
test_output[3594] = '{32'h430f1412};
/*############ DEBUG ############
test_input[28752:28759] = '{-5.44272983938, 18.1539221352, 22.7811982152, -94.8637424785, -43.2308322882, 99.8475605012, 72.7398897446, 85.6882179906};
test_label[3594] = '{-43.2308322882};
test_output[3594] = '{143.078393498};
############ END DEBUG ############*/
test_input[28760:28767] = '{32'hc2698ef5, 32'h42a20baa, 32'hc2954443, 32'h42657aff, 32'h41584d8c, 32'hc1227a21, 32'hc283d0b6, 32'hc2bdbe25};
test_label[3595] = '{32'hc283d0b6};
test_output[3595] = '{32'h4312ee30};
/*############ DEBUG ############
test_input[28760:28767] = '{-58.3896079944, 81.0227824507, -74.6333228299, 57.3701125304, 13.5189318911, -10.1548165094, -65.9076384765, -94.8713768086};
test_label[3595] = '{-65.9076384765};
test_output[3595] = '{146.930420927};
############ END DEBUG ############*/
test_input[28768:28775] = '{32'h426a0487, 32'h423312c4, 32'h42ab81e4, 32'hc22e376f, 32'hc2ba07d5, 32'h42a32d95, 32'h42615d43, 32'hc1c4c649};
test_label[3596] = '{32'hc2ba07d5};
test_output[3596] = '{32'h4332c8cf};
/*############ DEBUG ############
test_input[28768:28775] = '{58.5044213176, 44.7683241894, 85.7536957329, -43.5541359153, -93.0152956094, 81.5890253528, 56.3410754011, -24.5968180805};
test_label[3596] = '{-93.0152956094};
test_output[3596] = '{178.784406747};
############ END DEBUG ############*/
test_input[28776:28783] = '{32'hbfa7ebda, 32'hc28e52c2, 32'hc2c6025f, 32'hc27c419d, 32'hc204941f, 32'h42c4e256, 32'h4202e287, 32'hbfb53412};
test_label[3597] = '{32'hc2c6025f};
test_output[3597] = '{32'h4345725a};
/*############ DEBUG ############
test_input[28776:28783] = '{-1.31188512269, -71.1616358175, -99.0046274218, -63.0640767401, -33.1446512092, 98.4420646587, 32.7212170471, -1.41565155078};
test_label[3597] = '{-99.0046274218};
test_output[3597] = '{197.446692081};
############ END DEBUG ############*/
test_input[28784:28791] = '{32'h427da3fe, 32'hc29392b4, 32'hc1ad25db, 32'hc256cba3, 32'h42bd64be, 32'h42a0c825, 32'h4038df10, 32'hc27812c1};
test_label[3598] = '{32'h42bd64be};
test_output[3598] = '{32'h352464f5};
/*############ DEBUG ############
test_input[28784:28791] = '{63.4101497043, -73.786529408, -21.6434849765, -53.6988654751, 94.6967596021, 80.3909070443, 2.88861474474, -62.0183151758};
test_label[3598] = '{94.6967596021};
test_output[3598] = '{6.12416750322e-07};
############ END DEBUG ############*/
test_input[28792:28799] = '{32'h423fd0ac, 32'hc2a122fc, 32'hc24c962e, 32'hc2c318c0, 32'h425935aa, 32'hc1a91bc4, 32'h42c567c3, 32'h428322e3};
test_label[3599] = '{32'hc1a91bc4};
test_output[3599] = '{32'h42efaeb4};
/*############ DEBUG ############
test_input[28792:28799] = '{47.9537826467, -80.5683322476, -51.1466596634, -97.5483391881, 54.3024060474, -21.1385572766, 98.7026572672, 65.5681358472};
test_label[3599] = '{-21.1385572766};
test_output[3599] = '{119.841214544};
############ END DEBUG ############*/
test_input[28800:28807] = '{32'hc21a26a4, 32'h41a23373, 32'h42755887, 32'h4110c207, 32'hc1a8bf2b, 32'h41a654e0, 32'hc23acab8, 32'h42c1fcb3};
test_label[3600] = '{32'hc1a8bf2b};
test_output[3600] = '{32'h42ec2c7e};
/*############ DEBUG ############
test_input[28800:28807] = '{-38.5377334512, 20.2751226153, 61.3364522129, 9.04736952365, -21.0933431349, 20.7914433268, -46.6979677191, 96.993556212};
test_label[3600] = '{-21.0933431349};
test_output[3600] = '{118.086899347};
############ END DEBUG ############*/
test_input[28808:28815] = '{32'hc29c6658, 32'hc23b85a1, 32'hc23e0f7b, 32'hc2c1ebd2, 32'hc1d9d4c7, 32'hc2a6dbce, 32'hc1d1d5b1, 32'h4205e2c2};
test_label[3601] = '{32'hc29c6658};
test_output[3601] = '{32'h42df57b9};
/*############ DEBUG ############
test_input[28808:28815] = '{-78.1998889131, -46.8804972216, -47.5151187351, -96.960589026, -27.2288957506, -83.4293026724, -26.2293422012, 33.4714442334};
test_label[3601] = '{-78.1998889131};
test_output[3601] = '{111.671333146};
############ END DEBUG ############*/
test_input[28816:28823] = '{32'h429eb201, 32'hc1027f5e, 32'hc191030c, 32'hc2a2b83c, 32'h42899fe2, 32'h4282bc94, 32'h424efba3, 32'h4257702a};
test_label[3602] = '{32'h429eb201};
test_output[3602] = '{32'h37e613e2};
/*############ DEBUG ############
test_input[28816:28823] = '{79.3476640838, -8.1560958449, -18.1264885861, -81.3598357309, 68.812270538, 65.3683148759, 51.7457391703, 53.8595361328};
test_label[3602] = '{79.3476640838};
test_output[3602] = '{2.74273949688e-05};
############ END DEBUG ############*/
test_input[28824:28831] = '{32'h428934d7, 32'hc074cfa7, 32'h42bc80a5, 32'hc2b0fe73, 32'hc24e04fe, 32'hc2393e3b, 32'h42307b02, 32'h41ebcef7};
test_label[3603] = '{32'h42307b02};
test_output[3603] = '{32'h42488647};
/*############ DEBUG ############
test_input[28824:28831] = '{68.6032058398, -3.82517412564, 94.2512555555, -88.4969739507, -51.5048750075, -46.3107709519, 44.1201262115, 29.4760561274};
test_label[3603] = '{44.1201262115};
test_output[3603] = '{50.131129344};
############ END DEBUG ############*/
test_input[28832:28839] = '{32'hc28a87e7, 32'h4291f05b, 32'hc2a608bc, 32'h42a138b0, 32'hc2b2600e, 32'h42b055f6, 32'h41d6f134, 32'hc24bd15c};
test_label[3604] = '{32'hc24bd15c};
test_output[3604] = '{32'h430b1f74};
/*############ DEBUG ############
test_input[28832:28839] = '{-69.2654369653, 72.9694444996, -83.0170575165, 80.6107159086, -89.1876069199, 88.1678896574, 26.8677742401, -50.9544534158};
test_label[3604] = '{-50.9544534158};
test_output[3604] = '{139.122865537};
############ END DEBUG ############*/
test_input[28840:28847] = '{32'hc296de14, 32'hc2b3162e, 32'h423bf85c, 32'hc29fa775, 32'h42b22a05, 32'h42b9830b, 32'h4298afdc, 32'hc28a909a};
test_label[3605] = '{32'h42b22a05};
test_output[3605] = '{32'h406cbb67};
/*############ DEBUG ############
test_input[28840:28847] = '{-75.4337454893, -89.5433196447, 46.9925382889, -79.8270641384, 89.0820673674, 92.7559442139, 76.343478185, -69.2824243724};
test_label[3605] = '{89.0820673674};
test_output[3605] = '{3.69893813969};
############ END DEBUG ############*/
test_input[28848:28855] = '{32'hc27cd005, 32'hc206b93a, 32'hc0cdbfaa, 32'hc1237d57, 32'h42811f3e, 32'hc016d4aa, 32'h42855670, 32'h42c67e6d};
test_label[3606] = '{32'hc206b93a};
test_output[3606] = '{32'h4304ed85};
/*############ DEBUG ############
test_input[28848:28855] = '{-63.203144545, -33.6808867986, -6.42964658192, -10.2181004653, 64.5610172793, -2.35672988104, 66.6688221286, 99.2469241742};
test_label[3606] = '{-33.6808867986};
test_output[3606] = '{132.927810973};
############ END DEBUG ############*/
test_input[28856:28863] = '{32'hc271f146, 32'hc292e2aa, 32'hc29fc927, 32'hc1a056cd, 32'hc1a96f9f, 32'h42a8f202, 32'hc1c1962e, 32'hc281fca3};
test_label[3607] = '{32'hc1a056cd};
test_output[3607] = '{32'h42d107b6};
/*############ DEBUG ############
test_input[28856:28863] = '{-60.4856192184, -73.4427015517, -79.8928761912, -20.0423835891, -21.1795033733, 84.4726733555, -24.1983295815, -64.9934282076};
test_label[3607] = '{-20.0423835891};
test_output[3607] = '{104.515056945};
############ END DEBUG ############*/
test_input[28864:28871] = '{32'h427b95bd, 32'hc2c2cdd2, 32'h42c74759, 32'h424e9b2b, 32'hc2b17a97, 32'hc2935b0d, 32'hc1fd63bd, 32'hc1c1ceba};
test_label[3608] = '{32'h427b95bd};
test_output[3608] = '{32'h4212f8f6};
/*############ DEBUG ############
test_input[28864:28871] = '{62.8962294706, -97.4019933657, 99.6393543893, 51.6515316026, -88.7394306714, -73.6778356121, -31.6737012356, -24.2259408915};
test_label[3608] = '{62.8962294706};
test_output[3608] = '{36.7431249187};
############ END DEBUG ############*/
test_input[28872:28879] = '{32'h42395970, 32'h407379ae, 32'hc1dc6985, 32'hc1b18a0b, 32'h413fc6e2, 32'hc2ac7713, 32'hc26d1ab9, 32'h4138925f};
test_label[3609] = '{32'h4138925f};
test_output[3609] = '{32'h420b34d8};
/*############ DEBUG ############
test_input[28872:28879] = '{46.3373404718, 3.80430185532, -27.5515229661, -22.1924046176, 11.9860557315, -86.2325694246, -59.2760981883, 11.535735153};
test_label[3609] = '{11.535735153};
test_output[3609] = '{34.8016053188};
############ END DEBUG ############*/
test_input[28880:28887] = '{32'hc29a98c6, 32'hc006859c, 32'hc29dc914, 32'hc090624b, 32'hc22a9ca0, 32'h42705d44, 32'hc0d648f0, 32'hc1fbed0b};
test_label[3610] = '{32'hc22a9ca0};
test_output[3610] = '{32'h42cd7cf2};
/*############ DEBUG ############
test_input[28880:28887] = '{-77.2983883634, -2.10190497449, -78.892729807, -4.51199868838, -42.6529527582, 60.0910790068, -6.69640352962, -31.4907436449};
test_label[3610] = '{-42.6529527582};
test_output[3610] = '{102.744031765};
############ END DEBUG ############*/
test_input[28888:28895] = '{32'h3fa6a770, 32'hc1e90dd7, 32'h42a9629b, 32'hc229ed1d, 32'h42697ab2, 32'hc2a1bf69, 32'hc2411d5e, 32'h422bf54c};
test_label[3611] = '{32'h42697ab2};
test_output[3611] = '{32'h41d2950a};
/*############ DEBUG ############
test_input[28888:28895] = '{1.30198476282, -29.1317580784, 84.6925912622, -42.4815540594, 58.3698188516, -80.8738488824, -48.2786798141, 42.9895458394};
test_label[3611] = '{58.3698188516};
test_output[3611] = '{26.3227724107};
############ END DEBUG ############*/
test_input[28896:28903] = '{32'hc24c89d4, 32'hc1ab43ab, 32'hc15fcb27, 32'hc2c4d978, 32'h426a8be3, 32'h4136ad6f, 32'hc2724375, 32'hc2c2e706};
test_label[3612] = '{32'hc1ab43ab};
test_output[3612] = '{32'h42a016dc};
/*############ DEBUG ############
test_input[28896:28903] = '{-51.134598239, -21.408040229, -13.9870978556, -98.424740318, 58.6366096911, 11.4173420649, -60.5658760771, -97.4512200085};
test_label[3612] = '{-21.408040229};
test_output[3612] = '{80.04464992};
############ END DEBUG ############*/
test_input[28904:28911] = '{32'hc2b5b075, 32'hc2837349, 32'hc2a0a94d, 32'hc173f977, 32'h428192ae, 32'h42c460c2, 32'hc2c69a02, 32'hc2547e01};
test_label[3613] = '{32'h42c460c2};
test_output[3613] = '{32'h27600000};
/*############ DEBUG ############
test_input[28904:28911] = '{-90.8446400011, -65.7251667554, -80.3306629392, -15.2484044261, 64.7864872249, 98.1889791285, -99.3007932481, -53.1230506322};
test_label[3613] = '{98.1889791285};
test_output[3613] = '{3.10862446895e-15};
############ END DEBUG ############*/
test_input[28912:28919] = '{32'hc206facd, 32'hc2ae18b9, 32'hc2863092, 32'h41f31cd6, 32'h42b85196, 32'h41d904eb, 32'h4290ae73, 32'hc22502e5};
test_label[3614] = '{32'h41d904eb};
test_output[3614] = '{32'h4282105c};
/*############ DEBUG ############
test_input[28912:28919] = '{-33.7449217323, -87.0482877694, -67.0948646498, 30.3890802625, 92.1593493607, 27.127401015, 72.3407187712, -41.2528277037};
test_label[3614] = '{27.127401015};
test_output[3614] = '{65.0319483483};
############ END DEBUG ############*/
test_input[28920:28927] = '{32'hc2a04e70, 32'h41b8cbed, 32'h3fb0e8d7, 32'hc28546e4, 32'hc288c44b, 32'hc2b6cc39, 32'h42ab5679, 32'hc29c2956};
test_label[3615] = '{32'hc28546e4};
test_output[3615] = '{32'h43184eaf};
/*############ DEBUG ############
test_input[28920:28927] = '{-80.1532002574, 23.0995724116, 1.38210570469, -66.6384580163, -68.3833882417, -91.3988713672, 85.6688929127, -78.0807328262};
test_label[3615] = '{-66.6384580163};
test_output[3615] = '{152.307350929};
############ END DEBUG ############*/
test_input[28928:28935] = '{32'h4218d093, 32'h42c4e86c, 32'hc24082db, 32'hc256a602, 32'h42aa1844, 32'h42413348, 32'h41e1e5e9, 32'hc2b26243};
test_label[3616] = '{32'h41e1e5e9};
test_output[3616] = '{32'h428c6ef2};
/*############ DEBUG ############
test_input[28928:28935] = '{38.2036854094, 98.4539491665, -48.1277880713, -53.6621182722, 85.0473924626, 48.3000777239, 28.237260886, -89.1919179738};
test_label[3616] = '{28.237260886};
test_output[3616] = '{70.2166897857};
############ END DEBUG ############*/
test_input[28936:28943] = '{32'h412cbbbb, 32'hc2449b92, 32'hc1370f44, 32'hc1034ed2, 32'hc0dda483, 32'hc229299d, 32'hc29fa2c8, 32'h40c5f1c9};
test_label[3617] = '{32'hc0dda483};
test_output[3617] = '{32'h418ddb46};
/*############ DEBUG ############
test_input[28936:28943] = '{10.7958326548, -49.1519255664, -11.4412273969, -8.20674276672, -6.92633194629, -42.2906365299, -79.8179318799, 6.18576483654};
test_label[3617] = '{-6.92633194629};
test_output[3617] = '{17.7320665836};
############ END DEBUG ############*/
test_input[28944:28951] = '{32'hc27bcba4, 32'hc21d740c, 32'hc28b71bd, 32'hc155031d, 32'hc28555ab, 32'h4219e181, 32'hc1de4cee, 32'hc25f9c56};
test_label[3618] = '{32'hc27bcba4};
test_output[3618] = '{32'h42cad693};
/*############ DEBUG ############
test_input[28944:28951] = '{-62.9488682561, -39.3633265133, -69.7221484097, -13.3132601832, -66.6673192081, 38.4702190706, -27.7875628223, -55.9026724813};
test_label[3618] = '{-62.9488682561};
test_output[3618] = '{101.419087327};
############ END DEBUG ############*/
test_input[28952:28959] = '{32'hc2bf9377, 32'hc0853d10, 32'h429aacda, 32'h42991526, 32'hc29c815c, 32'h41617206, 32'hc21a82c9, 32'hc1b20e81};
test_label[3619] = '{32'hc2bf9377};
test_output[3619] = '{32'h432d7f74};
/*############ DEBUG ############
test_input[28952:28959] = '{-95.7880135721, -4.16370376051, 77.337597409, 76.5413060537, -78.2526512597, 14.090337559, -38.6277216554, -22.2570823616};
test_label[3619] = '{-95.7880135721};
test_output[3619] = '{173.497862893};
############ END DEBUG ############*/
test_input[28960:28967] = '{32'h42102151, 32'hc281d19e, 32'h427d4609, 32'h4160a891, 32'hc2216a5f, 32'hc21cfae7, 32'hc1afeb4c, 32'h414a87bd};
test_label[3620] = '{32'hc2216a5f};
test_output[3620] = '{32'h42cf5834};
/*############ DEBUG ############
test_input[28960:28967] = '{36.0325365584, -64.9094090625, 63.3183933019, 14.0411536337, -40.3538780871, -39.245020494, -21.9898907597, 12.6581395473};
test_label[3620] = '{-40.3538780871};
test_output[3620] = '{103.672271389};
############ END DEBUG ############*/
test_input[28968:28975] = '{32'hc060af17, 32'hc1b54cbe, 32'h421a48c8, 32'hc1de9b83, 32'hc2c62fa1, 32'h42a44806, 32'hc14d8d53, 32'h426f0bcd};
test_label[3621] = '{32'h421a48c8};
test_output[3621] = '{32'h422e4744};
/*############ DEBUG ############
test_input[28968:28975] = '{-3.51068660991, -22.6624724917, 38.5710739131, -27.8259326281, -99.093026419, 82.1406692876, -12.8470029287, 59.7615241807};
test_label[3621] = '{38.5710739131};
test_output[3621] = '{43.5695953747};
############ END DEBUG ############*/
test_input[28976:28983] = '{32'h41dcedef, 32'hc29f6e91, 32'h42c0d7a2, 32'hc20eb56f, 32'hc1942cd4, 32'h424262b3, 32'hc28d677e, 32'h42bde3ef};
test_label[3622] = '{32'h42bde3ef};
test_output[3622] = '{32'h3fd745b6};
/*############ DEBUG ############
test_input[28976:28983] = '{27.6161776392, -79.7159499958, 96.4211586624, -35.6771793693, -18.5218882006, 48.5963849146, -70.7021355939, 94.9451829115};
test_label[3622] = '{94.9451829115};
test_output[3622] = '{1.68181492522};
############ END DEBUG ############*/
test_input[28984:28991] = '{32'h41153222, 32'hc2a1badc, 32'hc213f8ae, 32'hc2c39d98, 32'hc254b295, 32'hc2c10b47, 32'hc174fc2e, 32'h411f9337};
test_label[3623] = '{32'hc254b295};
test_output[3623] = '{32'h427e45fb};
/*############ DEBUG ############
test_input[28984:28991] = '{9.32473978441, -80.8649633557, -36.9928516503, -97.8078007902, -53.1743979673, -96.5220245028, -15.3115677703, 9.97344119859};
test_label[3623] = '{-53.1743979673};
test_output[3623] = '{63.568340093};
############ END DEBUG ############*/
test_input[28992:28999] = '{32'hc2b8e15f, 32'hc2c2211b, 32'hc1f283d4, 32'hc27a50fd, 32'hc2a8f5e9, 32'hc2acdcc1, 32'hc28b9788, 32'h420f8363};
test_label[3624] = '{32'hc28b9788};
test_output[3624] = '{32'h42d3593a};
/*############ DEBUG ############
test_input[28992:28999] = '{-92.4401775143, -97.0646565685, -30.3143683886, -62.5790891895, -84.4802946672, -86.4311612842, -69.7959632398, 35.8783058343};
test_label[3624] = '{-69.7959632398};
test_output[3624] = '{105.674269074};
############ END DEBUG ############*/
test_input[29000:29007] = '{32'hc1d18ff9, 32'hc2998c61, 32'h42b8357d, 32'hc28a4b25, 32'hc28e3cf6, 32'hc2a5a555, 32'h418c2916, 32'h41ba4371};
test_label[3625] = '{32'hc2998c61};
test_output[3625] = '{32'h4328e0ef};
/*############ DEBUG ############
test_input[29000:29007] = '{-26.1952999333, -76.7741762421, 92.1044674359, -69.1467655002, -71.1190660114, -82.8229139302, 17.5200610806, 23.2829307788};
test_label[3625] = '{-76.7741762421};
test_output[3625] = '{168.878643678};
############ END DEBUG ############*/
test_input[29008:29015] = '{32'h429fd80f, 32'hc1da9329, 32'h4297b2f0, 32'h4261d4db, 32'hc11f3e45, 32'hc0f42295, 32'h3f421941, 32'hc0e05af2};
test_label[3626] = '{32'h3f421941};
test_output[3626] = '{32'h429e5c82};
/*############ DEBUG ############
test_input[29008:29015] = '{79.9219876351, -27.321856276, 75.8494892602, 56.4578652979, -9.95270269451, -7.62922140677, 0.758197821107, -7.01110155537};
test_label[3626] = '{0.758197821107};
test_output[3626] = '{79.1806811253};
############ END DEBUG ############*/
test_input[29016:29023] = '{32'h42b53280, 32'h42234437, 32'hc1dda974, 32'h41ef9a83, 32'hc24565ea, 32'hc1f9dc1a, 32'h41ec6cdb, 32'h42959c24};
test_label[3627] = '{32'hc1f9dc1a};
test_output[3627] = '{32'h42f3a986};
/*############ DEBUG ############
test_input[29016:29023] = '{90.5986311523, 40.8166161872, -27.7077403426, 29.9504450414, -49.3495247584, -31.2324719528, 29.5531529442, 74.8049604047};
test_label[3627] = '{-31.2324719528};
test_output[3627] = '{121.831103243};
############ END DEBUG ############*/
test_input[29024:29031] = '{32'hc2052917, 32'h42b012c4, 32'hc291b354, 32'h423807bb, 32'hc1b5ad9a, 32'hc257680a, 32'h41a1a9c6, 32'hc2758e3c};
test_label[3628] = '{32'hc1b5ad9a};
test_output[3628] = '{32'h42dd7e2a};
/*############ DEBUG ############
test_input[29024:29031] = '{-33.2901267483, 88.0366509642, -72.8502502288, 46.0075508964, -22.7097663154, -53.8516003728, 20.2078977876, -61.3889026631};
test_label[3628] = '{-22.7097663154};
test_output[3628] = '{110.74641728};
############ END DEBUG ############*/
test_input[29032:29039] = '{32'hc2a9ef91, 32'h42bd3be2, 32'hc12fb802, 32'h423ed337, 32'hc1909955, 32'hc1a6b644, 32'hc1cd3962, 32'hc298cfe9};
test_label[3629] = '{32'h42bd3be2};
test_output[3629] = '{32'h80000000};
/*############ DEBUG ############
test_input[29032:29039] = '{-84.9679017603, 94.6169581899, -10.9824241927, 47.7062639885, -18.0748694386, -20.8389959973, -25.6530185692, -76.4060762033};
test_label[3629] = '{94.6169581899};
test_output[3629] = '{-0.0};
############ END DEBUG ############*/
test_input[29040:29047] = '{32'hc1c232ae, 32'hc2b6ee16, 32'hc19b4bda, 32'hc23ebc36, 32'h427963c6, 32'h42a968d0, 32'hc22a0065, 32'hc28b6d8f};
test_label[3630] = '{32'hc23ebc36};
test_output[3630] = '{32'h43046375};
/*############ DEBUG ############
test_input[29040:29047] = '{-24.2747466518, -91.465008405, -19.4120377437, -47.6837979531, 62.3474358606, 84.7047096217, -42.5003838279, -69.7139822571};
test_label[3630] = '{-47.6837979531};
test_output[3630] = '{132.388507575};
############ END DEBUG ############*/
test_input[29048:29055] = '{32'h41b3be5a, 32'hc1b1d5bc, 32'h427f2667, 32'hc0c364a5, 32'hc28c61da, 32'hc280f35d, 32'hc20ecc58, 32'h40e952a3};
test_label[3631] = '{32'h427f2667};
test_output[3631] = '{32'h80000000};
/*############ DEBUG ############
test_input[29048:29055] = '{22.4679447067, -22.2293622091, 63.7875008342, -6.10603568748, -70.1911178374, -64.4753166513, -35.6995558216, 7.29133750251};
test_label[3631] = '{63.7875008342};
test_output[3631] = '{-0.0};
############ END DEBUG ############*/
test_input[29056:29063] = '{32'h42b71cf2, 32'hc2c4182f, 32'hc2b50256, 32'h4255ff17, 32'hc2b8c7c6, 32'hc0aaa572, 32'h4296d161, 32'h42a598e6};
test_label[3632] = '{32'hc2b8c7c6};
test_output[3632] = '{32'h4337f266};
/*############ DEBUG ############
test_input[29056:29063] = '{91.5565346955, -98.0472357078, -90.5045601867, 53.4991114628, -92.3901826971, -5.33269584873, 75.4089432278, 82.7986285587};
test_label[3632] = '{-92.3901826971};
test_output[3632] = '{183.946874691};
############ END DEBUG ############*/
test_input[29064:29071] = '{32'hc2781af3, 32'h42348d0d, 32'h424a77ce, 32'h415b74af, 32'h421b3992, 32'h424df79b, 32'h40a17a4d, 32'h41030c69};
test_label[3633] = '{32'h424a77ce};
test_output[3633] = '{32'h3f9cbd9c};
/*############ DEBUG ############
test_input[29064:29071] = '{-62.0263185866, 45.1377459974, 50.6169950786, 13.7159870985, 38.806222495, 51.491800377, 5.04617942163, 8.19053014095};
test_label[3633] = '{50.6169950786};
test_output[3633] = '{1.22453636565};
############ END DEBUG ############*/
test_input[29072:29079] = '{32'hc1eea73d, 32'hc2b6a14b, 32'hc29b0d14, 32'h420839da, 32'hc24e958b, 32'hc224cdee, 32'h428112cb, 32'hc222f267};
test_label[3634] = '{32'hc29b0d14};
test_output[3634] = '{32'h430e0fef};
/*############ DEBUG ############
test_input[29072:29079] = '{-29.8316590997, -91.3150284952, -77.525541784, 34.0564957958, -51.6460376021, -41.2011049133, 64.5367056712, -40.7367216185};
test_label[3634] = '{-77.525541784};
test_output[3634] = '{142.062247455};
############ END DEBUG ############*/
test_input[29080:29087] = '{32'hc2a812e8, 32'h42b274f6, 32'hc23f5a93, 32'h42964e7a, 32'h42bc3199, 32'hc2665ea4, 32'h42a0ad41, 32'hc2a93db0};
test_label[3635] = '{32'hc2a812e8};
test_output[3635] = '{32'h43322436};
/*############ DEBUG ############
test_input[29080:29087] = '{-84.036924326, 89.2284359205, -47.8384519784, 75.1532709096, 94.0968726757, -57.5924234977, 80.3383865029, -84.6204863825};
test_label[3635] = '{-84.036924326};
test_output[3635] = '{178.141454046};
############ END DEBUG ############*/
test_input[29088:29095] = '{32'h416180fb, 32'hc18a10f0, 32'hc2844d92, 32'hc1c7583c, 32'h4292484f, 32'h42c7616c, 32'hc2afe820, 32'h42bd8af9};
test_label[3636] = '{32'hc2844d92};
test_output[3636] = '{32'h4325d95c};
/*############ DEBUG ############
test_input[29088:29095] = '{14.0939892887, -17.258270073, -66.1515061387, -24.9180827278, 73.141226375, 99.6902754628, -87.9533728408, 94.7714289033};
test_label[3636] = '{-66.1515061387};
test_output[3636] = '{165.849062585};
############ END DEBUG ############*/
test_input[29096:29103] = '{32'hc2b05132, 32'h41c0f24d, 32'h42185275, 32'hc298942b, 32'h41c5e32e, 32'hc299cb4f, 32'h40ea90bf, 32'h41f467f3};
test_label[3637] = '{32'h41f467f3};
test_output[3637] = '{32'h40f0f84b};
/*############ DEBUG ############
test_input[29096:29103] = '{-88.1585861626, 24.1183111381, 38.0805257958, -76.2893895005, 24.7359274801, -76.8970886619, 7.33016931826, 30.5507557548};
test_label[3637] = '{30.5507557548};
test_output[3637] = '{7.53030922233};
############ END DEBUG ############*/
test_input[29104:29111] = '{32'hc28a27ee, 32'h415321c9, 32'h42a6d6ce, 32'hc265f89f, 32'h429d8ac0, 32'h42b9aa18, 32'hc231f589, 32'hc295a1d5};
test_label[3638] = '{32'hc265f89f};
test_output[3638] = '{32'h43165339};
/*############ DEBUG ############
test_input[29104:29111] = '{-69.0779845039, 13.1957485897, 83.4195440017, -57.4927944743, 78.7709988685, 92.8322164206, -44.489778981, -74.8160816899};
test_label[3638] = '{-57.4927944743};
test_output[3638] = '{150.325093356};
############ END DEBUG ############*/
test_input[29112:29119] = '{32'h424bd192, 32'hc25ee95c, 32'hc116dfbb, 32'h42c6aaca, 32'h41e2b821, 32'hc1f8eff3, 32'h4287a8b0, 32'hc2beaead};
test_label[3639] = '{32'h4287a8b0};
test_output[3639] = '{32'h41fc086a};
/*############ DEBUG ############
test_input[29112:29119] = '{50.9546569304, -55.7278913033, -9.42962168848, 99.3335751672, 28.3399069659, -31.117163626, 67.8294666829, -95.3411666905};
test_label[3639] = '{67.8294666829};
test_output[3639] = '{31.5041084843};
############ END DEBUG ############*/
test_input[29120:29127] = '{32'hc133fd52, 32'hc0c33437, 32'h41ca84be, 32'hc2aeeb86, 32'h417341a1, 32'h420cbac1, 32'hc228807f, 32'h425c2791};
test_label[3640] = '{32'hc133fd52};
test_output[3640] = '{32'h42849373};
/*############ DEBUG ############
test_input[29120:29127] = '{-11.2493460519, -6.10012408897, 25.3148155788, -87.4600041628, 15.2035227637, 35.1823768729, -42.1254840953, 55.0386403041};
test_label[3640] = '{-11.2493460519};
test_output[3640] = '{66.2879863583};
############ END DEBUG ############*/
test_input[29128:29135] = '{32'hc2363315, 32'hc1d221c4, 32'h42c486af, 32'h40874b53, 32'hc190ba3d, 32'hc188d6d4, 32'h410af387, 32'h41d3fb93};
test_label[3641] = '{32'hc1d221c4};
test_output[3641] = '{32'h42f90f20};
/*############ DEBUG ############
test_input[29128:29135] = '{-45.5498832449, -26.2664862827, 98.2630563058, 4.22794469695, -18.0909363123, -17.1048958411, 8.68445462903, 26.4978397916};
test_label[3641] = '{-26.2664862827};
test_output[3641] = '{124.529542588};
############ END DEBUG ############*/
test_input[29136:29143] = '{32'hc288c661, 32'hc279d646, 32'hc2220b77, 32'hc12a2a33, 32'hc1a95129, 32'h42827c4b, 32'h4209df55, 32'hc1a6a2aa};
test_label[3642] = '{32'hc12a2a33};
test_output[3642] = '{32'h4297c192};
/*############ DEBUG ############
test_input[29136:29143] = '{-68.3874567333, -62.4592497133, -40.5111946997, -10.6353025804, -21.164629476, 65.2427616966, 34.4680992433, -20.8294260141};
test_label[3642] = '{-10.6353025804};
test_output[3642] = '{75.878064277};
############ END DEBUG ############*/
test_input[29144:29151] = '{32'hc072f317, 32'h41f43096, 32'h41e53470, 32'hc25f6d07, 32'h429424ef, 32'hc26a4c5e, 32'h419170f8, 32'h41c0c751};
test_label[3643] = '{32'hc25f6d07};
test_output[3643] = '{32'h4301edb9};
/*############ DEBUG ############
test_input[29144:29151] = '{-3.79608690744, 30.5237240192, 28.6506050676, -55.8564714286, 74.0721338731, -58.5745760941, 18.1801612672, 24.0973234146};
test_label[3643] = '{-55.8564714286};
test_output[3643] = '{129.928605302};
############ END DEBUG ############*/
test_input[29152:29159] = '{32'hc211022c, 32'hc28f2095, 32'h42c47fef, 32'h42b18720, 32'h42975316, 32'h422622af, 32'h41c71f50, 32'hc24973db};
test_label[3644] = '{32'hc28f2095};
test_output[3644] = '{32'h4329d047};
/*############ DEBUG ############
test_input[29152:29159] = '{-36.2521210383, -71.5636368666, 98.2498740775, 88.7639197431, 75.6622754396, 41.5338715218, 24.8902896228, -50.3631393725};
test_label[3644] = '{-71.5636368666};
test_output[3644] = '{169.813586852};
############ END DEBUG ############*/
test_input[29160:29167] = '{32'h42b4856d, 32'hc2186099, 32'hc2758af1, 32'hc2013dc7, 32'hc115801e, 32'hc271ff9b, 32'hc2a652aa, 32'h426f9ea6};
test_label[3645] = '{32'hc271ff9b};
test_output[3645] = '{32'h4316c29d};
/*############ DEBUG ############
test_input[29160:29167] = '{90.2605993807, -38.0943335232, -61.3856847797, -32.3103285077, -9.34377877224, -60.4996137494, -83.1614543488, 59.9049293137};
test_label[3645] = '{-60.4996137494};
test_output[3645] = '{150.76021313};
############ END DEBUG ############*/
test_input[29168:29175] = '{32'hc190679e, 32'h429da9e1, 32'hc29eb629, 32'h41dcd6b5, 32'h4290218e, 32'hc2276ae2, 32'hc26e23de, 32'h3ff8c417};
test_label[3646] = '{32'h4290218e};
test_output[3646] = '{32'h40d88e9e};
/*############ DEBUG ############
test_input[29168:29175] = '{-18.0505939241, 78.8317983026, -79.3557847407, 27.6048375175, 72.0655400871, -41.8543781342, -59.5350247212, 1.94348416717};
test_label[3646] = '{72.0655400871};
test_output[3646] = '{6.76740954958};
############ END DEBUG ############*/
test_input[29176:29183] = '{32'h41a09c18, 32'h420ec421, 32'h4264bb37, 32'h429374fb, 32'h423658c5, 32'h424e0db3, 32'h422cd8cb, 32'h428c5dd4};
test_label[3647] = '{32'h424e0db3};
test_output[3647] = '{32'h41b1f2ce};
/*############ DEBUG ############
test_input[29176:29183] = '{20.0762185744, 35.6915318308, 57.1828268424, 73.7284795188, 45.5866891987, 51.5133769857, 43.2117118487, 70.1832554946};
test_label[3647] = '{51.5133769857};
test_output[3647] = '{22.2435560854};
############ END DEBUG ############*/
test_input[29184:29191] = '{32'h42b6088b, 32'hc29b85cf, 32'h427b960d, 32'hc0c3b6b8, 32'hbe74f22f, 32'hc19de69e, 32'hc2a7954e, 32'h428dc66e};
test_label[3648] = '{32'h42b6088b};
test_output[3648] = '{32'h30f90d0f};
/*############ DEBUG ############
test_input[29184:29191] = '{91.0166854632, -77.7613432505, 62.8965344825, -6.11605464736, -0.239205100008, -19.7376067327, -83.7916070634, 70.887559083};
test_label[3648] = '{91.0166854632};
test_output[3648] = '{1.81208459513e-09};
############ END DEBUG ############*/
test_input[29192:29199] = '{32'hc2497a1e, 32'hc2a4cec8, 32'h42ac7cb0, 32'hc1f91bba, 32'h42b5eb9b, 32'hc2891b9e, 32'h416c00d5, 32'h4288595a};
test_label[3649] = '{32'hc1f91bba};
test_output[3649] = '{32'h42f43719};
/*############ DEBUG ############
test_input[29192:29199] = '{-50.369254722, -82.4038705235, 86.2435305163, -31.138538977, 90.9601649993, -68.5539424152, 14.7502030722, 68.1745121352};
test_label[3649] = '{-31.138538977};
test_output[3649] = '{122.107609438};
############ END DEBUG ############*/
test_input[29200:29207] = '{32'hc28bc024, 32'h3fd0bfcb, 32'hc1af7e26, 32'hc2860bb3, 32'h428a4ef0, 32'h4154c732, 32'hc06c1175, 32'h4277597c};
test_label[3650] = '{32'h4154c732};
test_output[3650] = '{32'h425f6cc2};
/*############ DEBUG ############
test_input[29200:29207] = '{-69.8752766823, 1.63085311367, -21.9365964916, -67.0228535272, 69.1541774384, 13.2986316649, -3.68856544802, 61.8373865237};
test_label[3650] = '{13.2986316649};
test_output[3650] = '{55.8562098436};
############ END DEBUG ############*/
test_input[29208:29215] = '{32'hc2a1fc31, 32'h420d5cdf, 32'hc0a04ec9, 32'h4226e5bd, 32'h42599f18, 32'h4263f477, 32'hc1ce68a3, 32'h4268d24d};
test_label[3651] = '{32'hc2a1fc31};
test_output[3651] = '{32'h430b7979};
/*############ DEBUG ############
test_input[29208:29215] = '{-80.99256254, 35.3406960631, -5.00961721549, 41.724353915, 54.4053652786, 56.9887338416, -25.8010917493, 58.2053704307};
test_label[3651] = '{-80.99256254};
test_output[3651] = '{139.47450016};
############ END DEBUG ############*/
test_input[29216:29223] = '{32'hc28a330e, 32'hc2bbb7d8, 32'h4297b1af, 32'h4045d09f, 32'hc2c08345, 32'h41b8b794, 32'hc133652d, 32'h4120d894};
test_label[3652] = '{32'h4297b1af};
test_output[3652] = '{32'h80000000};
/*############ DEBUG ############
test_input[29216:29223] = '{-69.0997139733, -93.8590702878, 75.8470375587, 3.09085815696, -96.2563866831, 23.0896369556, -11.2122014105, 10.0528754888};
test_label[3652] = '{75.8470375587};
test_output[3652] = '{-0.0};
############ END DEBUG ############*/
test_input[29224:29231] = '{32'hc29ba4bc, 32'hc296f10d, 32'h42a755ed, 32'hc0480ff0, 32'hc2b34bef, 32'h42a0a29a, 32'h41f84352, 32'hc2c5bfa8};
test_label[3653] = '{32'hc29ba4bc};
test_output[3653] = '{32'h43218628};
/*############ DEBUG ############
test_input[29224:29231] = '{-77.821748402, -75.4708003775, 83.6678219602, -3.12597270521, -89.6483096875, 80.3175820476, 31.0328703308, -98.8743281371};
test_label[3653] = '{-77.821748402};
test_output[3653] = '{161.524045156};
############ END DEBUG ############*/
test_input[29232:29239] = '{32'h421c3ceb, 32'hc27d381e, 32'h42519c90, 32'hc2ae4809, 32'h42a40759, 32'h41fc8430, 32'h42c055d2, 32'hc26e527b};
test_label[3654] = '{32'h42519c90};
test_output[3654] = '{32'h422f0f14};
/*############ DEBUG ############
test_input[29232:29239] = '{39.0594885859, -63.3048007551, 52.4028918416, -87.1406930782, 82.0143482756, 31.5645453342, 96.1676141652, -59.580545541};
test_label[3654] = '{52.4028918416};
test_output[3654] = '{43.7647230369};
############ END DEBUG ############*/
test_input[29240:29247] = '{32'hc24cecff, 32'h42c0acc9, 32'h400bc597, 32'h42be30be, 32'hc1916e74, 32'h3f075158, 32'hc18b3fa5, 32'h429d385d};
test_label[3655] = '{32'h400bc597};
test_output[3655] = '{32'h42bcd07b};
/*############ DEBUG ############
test_input[29240:29247] = '{-51.2314412303, 96.3374679873, 2.18393485012, 95.0951974627, -18.1789321571, 0.528584936182, -17.4060765604, 78.6100872438};
test_label[3655] = '{2.18393485012};
test_output[3655] = '{94.4071887678};
############ END DEBUG ############*/
test_input[29248:29255] = '{32'h42aa2a2a, 32'hc28314e8, 32'h41f6c4fa, 32'hc22bf1fb, 32'h42b83521, 32'h4028532b, 32'h42aca916, 32'hc276921c};
test_label[3656] = '{32'hc22bf1fb};
test_output[3656] = '{32'h43071815};
/*############ DEBUG ############
test_input[29248:29255] = '{85.0823492204, -65.5408345664, 30.8461806108, -42.9863102524, 92.1037683508, 2.63007625145, 86.3302442373, -61.6426861989};
test_label[3656] = '{-42.9863102524};
test_output[3656] = '{135.09407196};
############ END DEBUG ############*/
test_input[29256:29263] = '{32'hc2a83f37, 32'h429a288b, 32'hc2b2de66, 32'hc26577e6, 32'hc253438d, 32'h426d0846, 32'hc28c0f11, 32'h401fc81f};
test_label[3657] = '{32'h426d0846};
test_output[3657] = '{32'h418e91a1};
/*############ DEBUG ############
test_input[29256:29263] = '{-84.1234649024, 77.0791867585, -89.4343708408, -57.3670896231, -52.815967168, 59.2580784808, -70.0294233839, 2.49658944756};
test_label[3657] = '{59.2580784808};
test_output[3657] = '{17.8211082959};
############ END DEBUG ############*/
test_input[29264:29271] = '{32'hc2a7caa8, 32'h414a33b1, 32'h422836ee, 32'h42c40d75, 32'h41f119a6, 32'h42884900, 32'hc1a17bfa, 32'hc18cb59d};
test_label[3658] = '{32'h42884900};
test_output[3658] = '{32'h41ef11d2};
/*############ DEBUG ############
test_input[29264:29271] = '{-83.8958113819, 12.637620059, 42.0536415026, 98.0262815566, 30.1375237216, 68.1425807233, -20.1855359298, -17.5886791373};
test_label[3658] = '{68.1425807233};
test_output[3658] = '{29.8837008333};
############ END DEBUG ############*/
test_input[29272:29279] = '{32'hc282b597, 32'hc2b21732, 32'h42064cfa, 32'hc1a57d36, 32'hc21e5fce, 32'h42861e29, 32'h42c5d7d5, 32'hc2b8a1d0};
test_label[3659] = '{32'hc21e5fce};
test_output[3659] = '{32'h430a83de};
/*############ DEBUG ############
test_input[29272:29279] = '{-65.3546645741, -89.0453030052, 33.5751727309, -20.686137792, -39.593559155, 67.0589080828, 98.9215446145, -92.3160392348};
test_label[3659] = '{-39.593559155};
test_output[3659] = '{138.515103769};
############ END DEBUG ############*/
test_input[29280:29287] = '{32'hbe845550, 32'h42365152, 32'h415d2528, 32'h4230ba19, 32'hc1111274, 32'h4258d075, 32'hc26e4a96, 32'hc23e7324};
test_label[3660] = '{32'h4230ba19};
test_output[3660] = '{32'h41205a5c};
/*############ DEBUG ############
test_input[29280:29287] = '{-0.258463376057, 45.5794141926, 13.8215715725, 44.1817358089, -9.06700517317, 54.2035721274, -59.5728392009, -47.6124433183};
test_label[3660] = '{44.1817358089};
test_output[3660] = '{10.0220604241};
############ END DEBUG ############*/
test_input[29288:29295] = '{32'h42ad27d7, 32'hc1925576, 32'hc11f4061, 32'h42465ba0, 32'h422ae6b8, 32'hc243b1c6, 32'hbfae0f15, 32'h42ac0140};
test_label[3661] = '{32'h42ac0140};
test_output[3661] = '{32'h3f82c59b};
/*############ DEBUG ############
test_input[29288:29295] = '{86.5778134516, -18.2917284091, -9.95321721793, 49.5894767836, 42.7253101729, -48.9236057277, -1.35983532435, 86.0024427809};
test_label[3661] = '{86.0024427809};
test_output[3661] = '{1.02165542403};
############ END DEBUG ############*/
test_input[29296:29303] = '{32'hc214d8ac, 32'h42549023, 32'h41ed67d3, 32'h428d4390, 32'hc23da528, 32'hc2aaace7, 32'hc28e1a2f, 32'h41bf7457};
test_label[3662] = '{32'hc28e1a2f};
test_output[3662] = '{32'h430daedf};
/*############ DEBUG ############
test_input[29296:29303] = '{-37.2115924195, 53.1407566856, 29.6756947573, 70.6319611594, -47.4112839814, -85.3376974591, -71.0511362233, 23.9318061198};
test_label[3662] = '{-71.0511362233};
test_output[3662] = '{141.683097408};
############ END DEBUG ############*/
test_input[29304:29311] = '{32'hc1f5aca1, 32'h41f7bf61, 32'hc2482f1e, 32'h429f511c, 32'h407d37f5, 32'h42930d55, 32'h41a8b73c, 32'h424dce53};
test_label[3663] = '{32'h41f7bf61};
test_output[3663] = '{32'h4242c4c1};
/*############ DEBUG ############
test_input[29304:29311] = '{-30.7092905773, 30.9684459971, -50.0460126223, 79.6584178241, 3.95654030048, 73.5260361604, 21.0894704151, 51.4514902014};
test_label[3663] = '{30.9684459971};
test_output[3663] = '{48.6921408761};
############ END DEBUG ############*/
test_input[29312:29319] = '{32'h4258c0a2, 32'hc29fa555, 32'h42224749, 32'h428de9ba, 32'hc2bca14b, 32'hc2a0fd14, 32'hc13ac7a2, 32'hc139e56c};
test_label[3664] = '{32'hc2bca14b};
test_output[3664] = '{32'h43254583};
/*############ DEBUG ############
test_input[29312:29319] = '{54.1881165619, -79.8229131484, 40.5696139554, 70.9565000932, -94.3150254424, -80.4942916712, -11.6737388149, -11.6185111669};
test_label[3664] = '{-94.3150254424};
test_output[3664] = '{165.271525588};
############ END DEBUG ############*/
test_input[29320:29327] = '{32'h42352dca, 32'h42a28029, 32'hc1314cd7, 32'h41eaa5ee, 32'h42794413, 32'hc23d2825, 32'hc011714a, 32'hc281e1eb};
test_label[3665] = '{32'h41eaa5ee};
test_output[3665] = '{32'h424fad5b};
/*############ DEBUG ############
test_input[29320:29327] = '{45.2947146127, 81.2503117511, -11.0812592642, 29.3310200251, 62.3164789025, -47.2892052261, -2.27253955265, -64.9412438143};
test_label[3665] = '{29.3310200251};
test_output[3665] = '{51.9192917319};
############ END DEBUG ############*/
test_input[29328:29335] = '{32'hc293fe6d, 32'hc17753a1, 32'hc14d618f, 32'hc286cf0b, 32'hc2b3da1c, 32'hc2151c9f, 32'hc235bf6f, 32'h3e182615};
test_label[3666] = '{32'hc14d618f};
test_output[3666] = '{32'h414fc22a};
/*############ DEBUG ############
test_input[29328:29335] = '{-73.9969270175, -15.4579174259, -12.8363178044, -67.4043783933, -89.9259965046, -37.2779505217, -45.4369486333, 0.148582764826};
test_label[3666] = '{-12.8363178044};
test_output[3666] = '{12.9849030307};
############ END DEBUG ############*/
test_input[29336:29343] = '{32'hc22ffd8f, 32'h423cb6d4, 32'h42a68516, 32'h4285ee4d, 32'hc1300db7, 32'h418bfd3e, 32'hc24675f9, 32'h4212e2d1};
test_label[3667] = '{32'h42a68516};
test_output[3667] = '{32'h33b404c4};
/*############ DEBUG ############
test_input[29336:29343] = '{-43.9976157563, 47.1785438259, 83.2599348291, 66.965432547, -11.0033479766, 17.4986538074, -49.6152062346, 36.721499363};
test_label[3667] = '{83.2599348291};
test_output[3667] = '{8.38277010748e-08};
############ END DEBUG ############*/
test_input[29344:29351] = '{32'h4186aeb8, 32'hc2987da5, 32'hc2aa01d8, 32'hc21bf320, 32'h42a7a9dc, 32'h4263e365, 32'h416000c7, 32'h426bd32f};
test_label[3668] = '{32'h4263e365};
test_output[3668] = '{32'h41d6e0a6};
/*############ DEBUG ############
test_input[29344:29351] = '{16.835311431, -76.24540108, -85.0036019851, -38.9874258412, 83.8317541944, 56.9720630995, 14.0001894195, 58.9562349157};
test_label[3668] = '{56.9720630995};
test_output[3668] = '{26.8596910949};
############ END DEBUG ############*/
test_input[29352:29359] = '{32'h414d13b9, 32'h4245abe2, 32'h41d19d05, 32'hc05b817f, 32'hc1dfa0ee, 32'h40a66483, 32'hc27aca59, 32'h42c7b366};
test_label[3669] = '{32'h4245abe2};
test_output[3669] = '{32'h4249bae9};
/*############ DEBUG ############
test_input[29352:29359] = '{12.817315098, 49.4178529226, 26.2016697609, -3.42977879238, -27.9535796021, 5.19976970633, -62.6976047911, 99.8503837668};
test_label[3669] = '{49.4178529226};
test_output[3669] = '{50.4325308442};
############ END DEBUG ############*/
test_input[29360:29367] = '{32'hc2a81a0e, 32'hc1878949, 32'h404b4000, 32'h42c0d0a3, 32'hc2a8b552, 32'h41bef5bf, 32'hc1fa596c, 32'h41f1bd31};
test_label[3670] = '{32'h41f1bd31};
test_output[3670] = '{32'h42846157};
/*############ DEBUG ############
test_input[29360:29367] = '{-84.050886277, -16.9420341496, 3.17578118299, 96.4074970651, -84.3541410743, 23.8699925017, -31.2936639556, 30.2173781425};
test_label[3670] = '{30.2173781425};
test_output[3670] = '{66.1901189226};
############ END DEBUG ############*/
test_input[29368:29375] = '{32'h42bf6e44, 32'hc1f39cda, 32'hc2865d4e, 32'hc281d6fa, 32'hc28f86a9, 32'h40426e9c, 32'h41913909, 32'h414e5e65};
test_label[3671] = '{32'hc2865d4e};
test_output[3671] = '{32'h4322e5c9};
/*############ DEBUG ############
test_input[29368:29375] = '{95.7153633756, -30.4515871429, -67.1822361105, -64.9198779662, -71.7630080717, 3.03800105044, 18.1528486492, 12.8980457687};
test_label[3671] = '{-67.1822361105};
test_output[3671] = '{162.897599486};
############ END DEBUG ############*/
test_input[29376:29383] = '{32'hc2b07a8b, 32'hc263fffc, 32'hc2a320e6, 32'hc2a5d59f, 32'hc2c590b5, 32'h4287e73e, 32'h423dbddf, 32'h42b4aa7b};
test_label[3672] = '{32'hc2c590b5};
test_output[3672] = '{32'h433d1d98};
/*############ DEBUG ############
test_input[29376:29383] = '{-88.2393420034, -56.9999863725, -81.5642556928, -82.9172317468, -98.7826338307, 67.951643791, 47.4354214881, 90.332971651};
test_label[3672] = '{-98.7826338307};
test_output[3672] = '{189.115605482};
############ END DEBUG ############*/
test_input[29384:29391] = '{32'h42c6f52d, 32'h41c81dab, 32'h42c4f64f, 32'h425391af, 32'hc2a29659, 32'hc1250a04, 32'h42aa8bf7, 32'h424234c1};
test_label[3673] = '{32'hc2a29659};
test_output[3673] = '{32'h4335161c};
/*############ DEBUG ############
test_input[29384:29391] = '{99.4788604918, 25.0144860933, 98.4810729351, 52.892271006, -81.293645839, -10.3149449248, 85.2733700551, 48.5515163251};
test_label[3673] = '{-81.293645839};
test_output[3673] = '{181.086364012};
############ END DEBUG ############*/
test_input[29392:29399] = '{32'h42740ca3, 32'hc2510e9a, 32'hc27645f6, 32'h3fcba73e, 32'hc2c4d8bd, 32'hc051f2f8, 32'hc2887102, 32'h42be2051};
test_label[3674] = '{32'hc2510e9a};
test_output[3674] = '{32'h431353cf};
/*############ DEBUG ############
test_input[29392:29399] = '{61.0123410667, -52.2642588342, -61.5683199223, 1.5910412911, -98.423314016, -3.2804545298, -68.220717023, 95.0631142079};
test_label[3674] = '{-52.2642588342};
test_output[3674] = '{147.327373042};
############ END DEBUG ############*/
test_input[29400:29407] = '{32'h40932a9d, 32'h42312946, 32'hc21dd10d, 32'h4179dd31, 32'h3f8675a0, 32'h41871cc6, 32'hc2933383, 32'h4228ea50};
test_label[3675] = '{32'hc21dd10d};
test_output[3675] = '{32'h42a7ba7f};
/*############ DEBUG ############
test_input[29400:29407] = '{4.59895199921, 44.2903065038, -39.4541501257, 15.6165018318, 1.05046459441, 16.8890493142, -73.600608584, 42.2288196034};
test_label[3675] = '{-39.4541501257};
test_output[3675] = '{83.8642506191};
############ END DEBUG ############*/
test_input[29408:29415] = '{32'h4285d3be, 32'h42993a83, 32'h4265c921, 32'hc21b0043, 32'h42b84d23, 32'h42b52c88, 32'h42a75333, 32'hc2bdd770};
test_label[3676] = '{32'hc21b0043};
test_output[3676] = '{32'h43031757};
/*############ DEBUG ############
test_input[29408:29415] = '{66.9135574083, 76.6142838861, 57.4464154887, -38.7502571372, 92.1506538609, 90.5869739075, 83.6625015553, -94.9207747947};
test_label[3676] = '{-38.7502571372};
test_output[3676] = '{131.091176149};
############ END DEBUG ############*/
test_input[29416:29423] = '{32'h42b04da8, 32'hc2aabcb6, 32'h41712718, 32'h427f3e7c, 32'hc2a309bc, 32'h42408a98, 32'hc2889fdf, 32'h4297b2ec};
test_label[3677] = '{32'hc2aabcb6};
test_output[3677] = '{32'h432d852f};
/*############ DEBUG ############
test_input[29416:29423] = '{88.1516759204, -85.3685740374, 15.0720448155, 63.8110181864, -81.5190121746, 48.1353456914, -68.3122488106, 75.8494575934};
test_label[3677] = '{-85.3685740374};
test_output[3677] = '{173.520254499};
############ END DEBUG ############*/
test_input[29424:29431] = '{32'hc19a504e, 32'h410ec3e9, 32'h42a885ea, 32'hbfc6d8a2, 32'h42c349b5, 32'hc14789ed, 32'hc2b2240f, 32'h421531c9};
test_label[3678] = '{32'hbfc6d8a2};
test_output[3678] = '{32'h42c66518};
/*############ DEBUG ############
test_input[29424:29431] = '{-19.2892115645, 8.92282990026, 84.2615509366, -1.55348605971, 97.643957331, -12.4711728618, -89.0704261678, 37.2986187503};
test_label[3678] = '{-1.55348605971};
test_output[3678] = '{99.1974449328};
############ END DEBUG ############*/
test_input[29432:29439] = '{32'hc20cd664, 32'h41fcceb5, 32'hc2bc9b73, 32'hc2a50cd8, 32'hc24c359f, 32'hc2a89be0, 32'h42848a30, 32'h42a0b14a};
test_label[3679] = '{32'h42a0b14a};
test_output[3679] = '{32'h354eccc2};
/*############ DEBUG ############
test_input[29432:29439] = '{-35.2093656408, 31.6009313009, -94.3036109313, -82.5250829726, -51.0523657002, -84.3044415939, 66.2698999566, 80.3462693115};
test_label[3679] = '{80.3462693115};
test_output[3679] = '{7.70389396486e-07};
############ END DEBUG ############*/
test_input[29440:29447] = '{32'h428954dc, 32'h41faa67e, 32'hc28f0f43, 32'hc12d3105, 32'hc288f121, 32'hc2bd6ae7, 32'hc28458ee, 32'h428905fe};
test_label[3680] = '{32'hc28458ee};
test_output[3680] = '{32'h43077562};
/*############ DEBUG ############
test_input[29440:29447] = '{68.6657438573, 31.3312958932, -71.5298112061, -10.8244679063, -68.4709552805, -94.7087930367, -66.173694225, 68.5117010021};
test_label[3680] = '{-66.173694225};
test_output[3680] = '{135.458527057};
############ END DEBUG ############*/
test_input[29448:29455] = '{32'h42ad3023, 32'h41de10ad, 32'h42b832c6, 32'hc1a17fe8, 32'hc21d1067, 32'h41790518, 32'h42b9a727, 32'h41ac5ab7};
test_label[3681] = '{32'h42b832c6};
test_output[3681] = '{32'h3f8fb8fa};
/*############ DEBUG ############
test_input[29448:29455] = '{86.5940170555, 27.7581428704, 92.0991685617, -20.187453281, -39.2660180285, 15.5637434712, 92.8264669217, 21.5442935826};
test_label[3681] = '{92.0991685617};
test_output[3681] = '{1.1228325379};
############ END DEBUG ############*/
test_input[29456:29463] = '{32'h418c0456, 32'hc29b72ce, 32'hc2427cab, 32'hc2b701e0, 32'h421bcf8f, 32'hc2bc9969, 32'hc180c6a4, 32'h42b990ff};
test_label[3682] = '{32'hc29b72ce};
test_output[3682] = '{32'h432a81e6};
/*############ DEBUG ############
test_input[29456:29463] = '{17.5021174435, -77.7242281681, -48.6217456309, -91.503664375, 38.9526936683, -94.2996281398, -16.0969927147, 92.7831936438};
test_label[3682] = '{-77.7242281681};
test_output[3682] = '{170.507421812};
############ END DEBUG ############*/
test_input[29464:29471] = '{32'hc25d40d9, 32'h40a4c528, 32'h41c83ae8, 32'h4234a77a, 32'h429a936f, 32'hc2452ba6, 32'hc21de595, 32'h423bea65};
test_label[3683] = '{32'hc25d40d9};
test_output[3683] = '{32'h430499ee};
/*############ DEBUG ############
test_input[29464:29471] = '{-55.313329655, 5.14906680657, 25.0287621031, 45.1635526683, 77.2879598733, -49.2926246722, -39.4742021983, 46.9789009965};
test_label[3683] = '{-55.313329655};
test_output[3683] = '{132.601289528};
############ END DEBUG ############*/
test_input[29472:29479] = '{32'hc2380b47, 32'h4216f862, 32'h42b965af, 32'h429ee922, 32'hc211c818, 32'hc26ba354, 32'hc28fafac, 32'hc290e88b};
test_label[3684] = '{32'hc211c818};
test_output[3684] = '{32'h430124de};
/*############ DEBUG ############
test_input[29472:29479] = '{-46.0110141705, 37.7425611583, 92.6986007921, 79.4553406275, -36.4454054364, -58.9095017805, -71.8431068344, -72.4541827233};
test_label[3684] = '{-36.4454054364};
test_output[3684] = '{129.144008001};
############ END DEBUG ############*/
test_input[29480:29487] = '{32'h42a01902, 32'hc00892af, 32'h421240ba, 32'hc255858f, 32'hc2795f61, 32'hc2937f59, 32'h425e2cc0, 32'hc26fced1};
test_label[3685] = '{32'hc255858f};
test_output[3685] = '{32'h43056de5};
/*############ DEBUG ############
test_input[29480:29487] = '{80.0488401023, -2.13395282748, 36.5632092625, -53.3804289473, -62.3431422567, -73.7487243354, 55.5437008352, -59.9519704979};
test_label[3685] = '{-53.3804289473};
test_output[3685] = '{133.42926905};
############ END DEBUG ############*/
test_input[29488:29495] = '{32'h428f8a24, 32'h42a135b8, 32'hc26fe285, 32'h42402eb4, 32'h4296ba72, 32'h41033b5c, 32'h41cc922d, 32'hc2bbfe24};
test_label[3686] = '{32'h42a135b8};
test_output[3686] = '{32'h3bb1d49d};
/*############ DEBUG ############
test_input[29488:29495] = '{71.7698078065, 80.6049200811, -59.9712114967, 48.0456075276, 75.3641500308, 8.20199199811, 25.5713750598, -93.9963653206};
test_label[3686] = '{80.6049200811};
test_output[3686] = '{0.00542695667093};
############ END DEBUG ############*/
test_input[29496:29503] = '{32'hc2b10a16, 32'hc20e5850, 32'hc274e9a1, 32'hc23f9d5b, 32'h42bce077, 32'hc2a8da7c, 32'hc1c7cd67, 32'h42a32b83};
test_label[3687] = '{32'h42bce077};
test_output[3687] = '{32'h362fa27e};
/*############ DEBUG ############
test_input[29496:29503] = '{-88.5197027401, -35.5862409644, -61.2281547273, -47.9036683223, 94.4384052412, -84.4267255995, -24.9752936861, 81.5849863377};
test_label[3687] = '{94.4384052412};
test_output[3687] = '{2.61716153222e-06};
############ END DEBUG ############*/
test_input[29504:29511] = '{32'h4286004a, 32'h41fdb970, 32'h427b9295, 32'h42a0305c, 32'h424610b8, 32'hc11bb13c, 32'h42409608, 32'h42bf1421};
test_label[3688] = '{32'h4286004a};
test_output[3688] = '{32'h41e44f5f};
/*############ DEBUG ############
test_input[29504:29511] = '{67.0005616756, 31.7155461297, 62.8931477079, 80.0944549198, 49.5163281294, -9.73077009706, 48.1465137272, 95.5393168879};
test_label[3688] = '{67.0005616756};
test_output[3688] = '{28.5387554084};
############ END DEBUG ############*/
test_input[29512:29519] = '{32'h4274be51, 32'hc229a35c, 32'h42a618cf, 32'hc22c78ce, 32'hc1bf4670, 32'h42938a70, 32'h42b19713, 32'h427ac005};
test_label[3689] = '{32'h4274be51};
test_output[3689] = '{32'h41dce631};
/*############ DEBUG ############
test_input[29512:29519] = '{61.1858561916, -42.409530841, 83.0484571167, -43.117972098, -23.9093926262, 73.7703892133, 88.7950662926, 62.6875206495};
test_label[3689] = '{61.1858561916};
test_output[3689] = '{27.6123989012};
############ END DEBUG ############*/
test_input[29520:29527] = '{32'hc2848f62, 32'h42b9f43c, 32'hc26339ea, 32'hc25d2b6c, 32'h4291a187, 32'h411ba8d5, 32'h42a43313, 32'hc20f4a7b};
test_label[3690] = '{32'hc25d2b6c};
test_output[3690] = '{32'h431444fa};
/*############ DEBUG ############
test_input[29520:29527] = '{-66.2800460166, 92.9770185228, -56.8065568382, -55.2924037019, 72.815480439, 9.72871866589, 82.0997569532, -35.8227339253};
test_label[3690] = '{-55.2924037019};
test_output[3690] = '{148.269441109};
############ END DEBUG ############*/
test_input[29528:29535] = '{32'hc1f3e94f, 32'h42830d55, 32'h41f8ab81, 32'hc0c2ad71, 32'h427494ce, 32'h4006819d, 32'h42960136, 32'hc2800284};
test_label[3691] = '{32'h427494ce};
test_output[3691] = '{32'h415db6c9};
/*############ DEBUG ############
test_input[29528:29535] = '{-30.4889206786, 65.5260388152, 31.0837420778, -6.08367225235, 61.1453188388, 2.10166104965, 75.0023668421, -64.0049137868};
test_label[3691] = '{61.1453188388};
test_output[3691] = '{13.8571256045};
############ END DEBUG ############*/
test_input[29536:29543] = '{32'hc2057996, 32'h408c404d, 32'h4135de77, 32'h42bd63db, 32'hc1727165, 32'hc29f5ee9, 32'hc29aafa9, 32'hc295e217};
test_label[3692] = '{32'h4135de77};
test_output[3692] = '{32'h42a6a80c};
/*############ DEBUG ############
test_input[29536:29543] = '{-33.3687365312, 4.38284920663, 11.3668124533, 94.6950312671, -15.1526839554, -79.6853709948, -77.3430883235, -74.9415847562};
test_label[3692] = '{11.3668124533};
test_output[3692] = '{83.3282188138};
############ END DEBUG ############*/
test_input[29544:29551] = '{32'hc2abda95, 32'hc2c42d58, 32'h428829e0, 32'hc20b970c, 32'hc21b74c8, 32'h422cf4d7, 32'h41d1d71b, 32'hc28ddbbc};
test_label[3693] = '{32'h41d1d71b};
test_output[3693] = '{32'h42276833};
/*############ DEBUG ############
test_input[29544:29551] = '{-85.9269153856, -98.0885647359, 68.0817891186, -34.8975080805, -38.8640447984, 43.2391012935, 26.230031759, -70.929170036};
test_label[3693] = '{26.230031759};
test_output[3693] = '{41.8517573596};
############ END DEBUG ############*/
test_input[29552:29559] = '{32'h41c466ee, 32'h3f346b8b, 32'h41501210, 32'h421986df, 32'h42144290, 32'h41f45725, 32'h40e181ee, 32'h41c0efe7};
test_label[3694] = '{32'h41501210};
test_output[3694] = '{32'h41cceba9};
/*############ DEBUG ############
test_input[29552:29559] = '{24.5502588773, 0.70476599835, 13.0044093461, 38.3817116129, 37.0650035857, 30.5425513911, 7.04711064451, 24.1171402396};
test_label[3694] = '{13.0044093461};
test_output[3694] = '{25.6150678141};
############ END DEBUG ############*/
test_input[29560:29567] = '{32'hc1cc0c98, 32'h4213b50d, 32'h418fa72c, 32'hc24f747f, 32'h429ae86e, 32'hc268afd6, 32'h4106b5d8, 32'h425425cb};
test_label[3695] = '{32'h418fa72c};
test_output[3695] = '{32'h426dfd47};
/*############ DEBUG ############
test_input[29560:29567] = '{-25.5061495347, 36.926808556, 17.9566266939, -51.8637665899, 77.4539672112, -58.1717147439, 8.41939556803, 53.036906937};
test_label[3695] = '{17.9566266939};
test_output[3695] = '{59.4973405174};
############ END DEBUG ############*/
test_input[29568:29575] = '{32'hc2b9e345, 32'h42c7ee74, 32'hc1fb6b2c, 32'h41904aa0, 32'hc28445aa, 32'hc2932073, 32'hc24161a8, 32'hc14ee94e};
test_label[3696] = '{32'hc14ee94e};
test_output[3696] = '{32'h42e1cb9e};
/*############ DEBUG ############
test_input[29568:29575] = '{-92.9438827804, 99.9657275952, -31.4273297597, 18.0364373281, -66.1360661319, -73.5633741052, -48.3453670076, -12.9319593269};
test_label[3696] = '{-12.9319593269};
test_output[3696] = '{112.897686922};
############ END DEBUG ############*/
test_input[29576:29583] = '{32'h418cd3f8, 32'h4223255a, 32'hc2ae6922, 32'h42b51328, 32'h40963d4e, 32'h41e8508b, 32'h42a30449, 32'hc0c5b610};
test_label[3697] = '{32'h42a30449};
test_output[3697] = '{32'h41107775};
/*############ DEBUG ############
test_input[29576:29583] = '{17.6035010033, 40.7864769202, -87.20533786, 90.5374158692, 4.69498350852, 29.0393284962, 81.5083714881, -6.1784743233};
test_label[3697] = '{81.5083714881};
test_output[3697] = '{9.02916425096};
############ END DEBUG ############*/
test_input[29584:29591] = '{32'hc2a3dff6, 32'hc17ab39c, 32'h421926a7, 32'h42285628, 32'h41cb83cb, 32'h42b3e247, 32'hc2b6dd6a, 32'hc280174c};
test_label[3698] = '{32'h42b3e247};
test_output[3698] = '{32'h80000000};
/*############ DEBUG ############
test_input[29584:29591] = '{-81.9374238751, -15.6688500745, 38.2877468185, 42.0841367351, 25.4393521558, 89.94195021, -91.4324519023, -64.0455016196};
test_label[3698] = '{89.94195021};
test_output[3698] = '{-0.0};
############ END DEBUG ############*/
test_input[29592:29599] = '{32'h3ff46e52, 32'hbd2fd10a, 32'hc11b3261, 32'h42862c62, 32'h41aeb943, 32'hc1841a7e, 32'h4149d5fb, 32'h41507f2e};
test_label[3699] = '{32'h4149d5fb};
test_output[3699] = '{32'h4259e344};
/*############ DEBUG ############
test_input[29592:29599] = '{1.90961674715, -0.0429239645209, -9.69979974656, 67.0866814793, 21.840459187, -16.5129350956, 12.6147416266, 13.0310500207};
test_label[3699] = '{12.6147416266};
test_output[3699] = '{54.4719398526};
############ END DEBUG ############*/
test_input[29600:29607] = '{32'h42b33f5c, 32'hc290f22a, 32'hc23e05dd, 32'hc27c5270, 32'hc28ba879, 32'hc1d25428, 32'hc2a1a0da, 32'h41b8dc42};
test_label[3700] = '{32'h41b8dc42};
test_output[3700] = '{32'h4285084c};
/*############ DEBUG ############
test_input[29600:29607] = '{89.6237504983, -72.4729731076, -47.5057262767, -63.0805043168, -69.8290459971, -26.2910913501, -80.8141657422, 23.1075475398};
test_label[3700] = '{23.1075475398};
test_output[3700] = '{66.5162029585};
############ END DEBUG ############*/
test_input[29608:29615] = '{32'h425c9976, 32'h41b5b5cb, 32'h4232533a, 32'h420d6f17, 32'h428b3246, 32'h428f8f3f, 32'h4299fa24, 32'h42b55385};
test_label[3701] = '{32'h428f8f3f};
test_output[3701] = '{32'h41971117};
/*############ DEBUG ############
test_input[29608:29615] = '{55.149865925, 22.7137667637, 44.5812740471, 35.3584870202, 69.5981932914, 71.7797781778, 76.9885548627, 90.6631207422};
test_label[3701] = '{71.7797781778};
test_output[3701] = '{18.8833437227};
############ END DEBUG ############*/
test_input[29616:29623] = '{32'h42b5da7d, 32'hc29660a3, 32'hc23681ee, 32'h4259e878, 32'hc28dd704, 32'h41c8e55f, 32'h42b615f6, 32'h40f8f755};
test_label[3702] = '{32'h40f8f755};
test_output[3702] = '{32'h42a7cc85};
/*############ DEBUG ############
test_input[29616:29623] = '{90.9267341829, -75.1887404179, -45.6268860583, 54.4770198016, -70.9199508538, 25.1119981027, 91.0428898617, 7.78019180195};
test_label[3702] = '{7.78019180195};
test_output[3702] = '{83.8994529714};
############ END DEBUG ############*/
test_input[29624:29631] = '{32'h421bb297, 32'hc1b5474e, 32'h421b1e73, 32'h4262971b, 32'h42240027, 32'hc207dbce, 32'hc2249f0a, 32'h42bcd23c};
test_label[3703] = '{32'h421bb297};
test_output[3703] = '{32'h425df1e2};
/*############ DEBUG ############
test_input[29624:29631] = '{38.9244033583, -22.6598168105, 38.7797338024, 56.6475653989, 41.0001493578, -33.9646536779, -41.1553120141, 94.4106152732};
test_label[3703] = '{38.9244033583};
test_output[3703] = '{55.4862119149};
############ END DEBUG ############*/
test_input[29632:29639] = '{32'hc293bfb0, 32'h42236365, 32'hc292cab2, 32'hc2b6d527, 32'h42bd69dc, 32'h4181484f, 32'hc2161cdb, 32'hc2703a50};
test_label[3704] = '{32'h42236365};
test_output[3704] = '{32'h42577052};
/*############ DEBUG ############
test_input[29632:29639] = '{-73.8743864266, 40.8470649378, -73.3958921418, -91.41631092, 94.7067540024, 16.1603060639, -37.5281778856, -60.0569439303};
test_label[3704] = '{40.8470649378};
test_output[3704] = '{53.8596890645};
############ END DEBUG ############*/
test_input[29640:29647] = '{32'h424651b2, 32'hc20a22c1, 32'h41931a80, 32'h418e5adf, 32'h41dd4ec2, 32'hc19e27ff, 32'hc1377458, 32'hc2067eb0};
test_label[3705] = '{32'hc19e27ff};
test_output[3705] = '{32'h428ab2d9};
/*############ DEBUG ############
test_input[29640:29647] = '{49.5797792494, -34.5339399753, 18.387939851, 17.7943697602, 27.6634565911, -19.7695299467, -11.4659040275, -33.6237176831};
test_label[3705] = '{-19.7695299467};
test_output[3705] = '{69.3493091964};
############ END DEBUG ############*/
test_input[29648:29655] = '{32'hc2387e69, 32'hc2b402f3, 32'hc2052d9a, 32'hc24b9394, 32'h418244a7, 32'h42bd9219, 32'hc2b310c9, 32'hc2b351f8};
test_label[3706] = '{32'hc2b402f3};
test_output[3706] = '{32'h4338ca86};
/*############ DEBUG ############
test_input[29648:29655] = '{-46.1234481641, -90.0057628874, -33.2945326255, -50.8941186673, 16.2835208599, 94.785346252, -89.5327840728, -89.6600955599};
test_label[3706] = '{-90.0057628874};
test_output[3706] = '{184.791109139};
############ END DEBUG ############*/
test_input[29656:29663] = '{32'h4298acdc, 32'h41934237, 32'h40aa801e, 32'h413ec1b2, 32'hc114662c, 32'hc1d43491, 32'h4206eee8, 32'h42b60919};
test_label[3707] = '{32'h413ec1b2};
test_output[3707] = '{32'h429e30e3};
/*############ DEBUG ############
test_input[29656:29663] = '{76.3376173478, 18.407332282, 5.32813935684, 11.9222891149, -9.2749442549, -26.5256666737, 33.7333082468, 91.0177717128};
test_label[3707] = '{11.9222891149};
test_output[3707] = '{79.0954830191};
############ END DEBUG ############*/
test_input[29664:29671] = '{32'h429b7532, 32'hc2b5a4a8, 32'h40155895, 32'h41a0ac60, 32'h423d16f4, 32'h42358ce9, 32'h42b67389, 32'hc239f974};
test_label[3708] = '{32'h41a0ac60};
test_output[3708] = '{32'h428e4871};
/*############ DEBUG ############
test_input[29664:29671] = '{77.7288992106, -90.821590967, 2.33353154652, 20.0841683698, 47.2724169142, 45.3876078798, 91.2256578534, -46.4936070051};
test_label[3708] = '{20.0841683698};
test_output[3708] = '{71.141490859};
############ END DEBUG ############*/
test_input[29672:29679] = '{32'h429b57fd, 32'h418b4a09, 32'h42607fd2, 32'h424cb313, 32'hc29158fc, 32'h4283bf04, 32'hc08996cc, 32'hc2451474};
test_label[3709] = '{32'hc08996cc};
test_output[3709] = '{32'h42a3f16b};
/*############ DEBUG ############
test_input[29672:29679] = '{77.6718520458, 17.4111493057, 56.1248262005, 51.1748778413, -72.673800129, 65.8730798995, -4.29965781629, -49.2699721598};
test_label[3709] = '{-4.29965781629};
test_output[3709] = '{81.9715173763};
############ END DEBUG ############*/
test_input[29680:29687] = '{32'h4234f8db, 32'hc1b1afa6, 32'h41fe6554, 32'hc229b642, 32'hc2b5172b, 32'hc26720a8, 32'h3e889a5e, 32'hc2884fb8};
test_label[3710] = '{32'h4234f8db};
test_output[3710] = '{32'h35c2b1a0};
/*############ DEBUG ############
test_input[29680:29687] = '{45.2430210494, -22.2107661299, 31.799476238, -42.427986143, -90.545248656, -57.7818908604, 0.26680271506, -68.1556992476};
test_label[3710] = '{45.2430210494};
test_output[3710] = '{1.45058224093e-06};
############ END DEBUG ############*/
test_input[29688:29695] = '{32'h42580af4, 32'h422227fa, 32'h428029c8, 32'hc21cca56, 32'h3f47c93b, 32'hc27e8138, 32'hc25ecb8a, 32'h4292b58d};
test_label[3711] = '{32'h428029c8};
test_output[3711] = '{32'h41145e85};
/*############ DEBUG ############
test_input[29688:29695] = '{54.0106968093, 40.5390406724, 64.0816065492, -39.1975923481, 0.78041431275, -63.6261886107, -55.6987683926, 73.3545883382};
test_label[3711] = '{64.0816065492};
test_output[3711] = '{9.27307571661};
############ END DEBUG ############*/
test_input[29696:29703] = '{32'h42ac5e93, 32'h4253d4e4, 32'hc1127aef, 32'hc1ca42ef, 32'h4292d0f2, 32'hc298dc55, 32'h411ef999, 32'h4048e87f};
test_label[3712] = '{32'hc298dc55};
test_output[3712] = '{32'h43229d74};
/*############ DEBUG ############
test_input[29696:29703] = '{86.1847163414, 52.95789987, -9.15501320706, -25.2826822997, 73.4080955382, -76.4303375987, 9.93593725944, 3.13919035968};
test_label[3712] = '{-76.4303375987};
test_output[3712] = '{162.615056766};
############ END DEBUG ############*/
test_input[29704:29711] = '{32'h414fa144, 32'h423bb1a0, 32'h41cae75c, 32'h423820b9, 32'h426de215, 32'h421c94f8, 32'h4265f81b, 32'h429e9c42};
test_label[3713] = '{32'h423bb1a0};
test_output[3713] = '{32'h420186e4};
/*############ DEBUG ############
test_input[29704:29711] = '{12.9768719128, 46.9234616501, 25.3629692945, 46.0319562559, 59.4707817749, 39.1454755475, 57.4922918886, 79.3051924519};
test_label[3713] = '{46.9234616501};
test_output[3713] = '{32.3817308046};
############ END DEBUG ############*/
test_input[29712:29719] = '{32'h428706ba, 32'hc249c964, 32'hc20d5402, 32'h4281679d, 32'hc2b368ce, 32'h4214247e, 32'hc2361d44, 32'hc17d0ec1};
test_label[3714] = '{32'h4214247e};
test_output[3714] = '{32'h41f44990};
/*############ DEBUG ############
test_input[29712:29719] = '{67.5131351117, -50.4466688074, -35.332039324, 64.7023662523, -89.7046996719, 37.0356352488, -45.5285813312, -15.8161023249};
test_label[3714] = '{37.0356352488};
test_output[3714] = '{30.5359184966};
############ END DEBUG ############*/
test_input[29720:29727] = '{32'hc295fb85, 32'hc2a5c31e, 32'hc2bf2dfb, 32'h42b7b30d, 32'h41d9588f, 32'hc173c57b, 32'hc2b64021, 32'hc25af1f8};
test_label[3715] = '{32'hc173c57b};
test_output[3715] = '{32'h42d62bbd};
/*############ DEBUG ############
test_input[29720:29727] = '{-74.9912470632, -82.8810914759, -95.5898048544, 91.8497120265, 27.1682421634, -15.2357130353, -91.1252528422, -54.7362979479};
test_label[3715] = '{-15.2357130353};
test_output[3715] = '{107.085425062};
############ END DEBUG ############*/
test_input[29728:29735] = '{32'hc125958d, 32'hc199969e, 32'h41cf34bc, 32'h42b14aad, 32'hc29151ab, 32'h40fac0af, 32'h42c2d0b3, 32'h42a5c96c};
test_label[3716] = '{32'h42a5c96c};
test_output[3716] = '{32'h41683ada};
/*############ DEBUG ############
test_input[29728:29735] = '{-10.349011748, -19.1985437491, 25.900748413, 88.6458501464, -72.6595041239, 7.83602071152, 97.4076133201, 82.8934020387};
test_label[3716] = '{82.8934020387};
test_output[3716] = '{14.5143683746};
############ END DEBUG ############*/
test_input[29736:29743] = '{32'hc2026ce7, 32'hc24e6b88, 32'h42577c93, 32'hc2b35515, 32'h426e88c3, 32'h425068ec, 32'hc06b40b3, 32'h419ea00f};
test_label[3717] = '{32'hc24e6b88};
test_output[3717] = '{32'h42de7c07};
/*############ DEBUG ############
test_input[29736:29743] = '{-32.6063488358, -51.6050105388, 53.8716561916, -89.6661761096, 59.6335569772, 52.10246341, -3.6758239126, 19.8281542088};
test_label[3717] = '{-51.6050105388};
test_output[3717] = '{111.242242036};
############ END DEBUG ############*/
test_input[29744:29751] = '{32'hc255ab35, 32'h426624b9, 32'h4187ebda, 32'hc2c6902b, 32'h4106abf9, 32'hc1685b8d, 32'h42139783, 32'hc2afde24};
test_label[3718] = '{32'h4106abf9};
test_output[3718] = '{32'h424479bb};
/*############ DEBUG ############
test_input[29744:29751] = '{-53.4171955187, 57.5358615437, 16.9901627379, -99.2815785733, 8.41698595713, -14.5223514362, 36.8979599791, -87.9338688438};
test_label[3718] = '{8.41698595713};
test_output[3718] = '{49.1188755876};
############ END DEBUG ############*/
test_input[29752:29759] = '{32'h425d5de3, 32'h429c5c55, 32'h4267f0b5, 32'hc28aba25, 32'h42947e20, 32'hc2a470c6, 32'hc1e16215, 32'hc2bc20d3};
test_label[3719] = '{32'h42947e20};
test_output[3719] = '{32'h407d0424};
/*############ DEBUG ############
test_input[29752:29759] = '{55.3416880187, 78.1803364696, 57.985067355, -69.3635604631, 74.2463351357, -82.2202605891, -28.1728912965, -94.0641068795};
test_label[3719] = '{74.2463351357};
test_output[3719] = '{3.95337762569};
############ END DEBUG ############*/
test_input[29760:29767] = '{32'hc2bb613a, 32'hc05da90b, 32'h418a765c, 32'h42383127, 32'hc19e2aaf, 32'hc2812ba5, 32'h41b2605f, 32'h42a45bf0};
test_label[3720] = '{32'h42a45bf0};
test_output[3720] = '{32'h25000000};
/*############ DEBUG ############
test_input[29760:29767] = '{-93.6898930499, -3.46344261168, 17.3077934903, 46.0480019888, -19.7708423366, -64.5852409848, 22.2970558702, 82.1795640947};
test_label[3720] = '{82.1795640947};
test_output[3720] = '{1.11022302463e-16};
############ END DEBUG ############*/
test_input[29768:29775] = '{32'hc2340137, 32'hc2c47492, 32'hc01853d7, 32'hc2973243, 32'hc22d203d, 32'hc2989e26, 32'h421e7605, 32'h4295bcfe};
test_label[3721] = '{32'hc2989e26};
test_output[3721] = '{32'h43172d92};
/*############ DEBUG ############
test_input[29768:29775] = '{-45.0011870328, -98.2276776009, -2.38011726581, -75.5981649655, -43.2814816789, -76.3088817592, 39.6152551097, 74.8691253999};
test_label[3721] = '{-76.3088817592};
test_output[3721] = '{151.178007159};
############ END DEBUG ############*/
test_input[29776:29783] = '{32'hc2c56860, 32'h427a696b, 32'hc265fd24, 32'hc1e76cc0, 32'h42a269c0, 32'hc08f0c64, 32'h408a05fa, 32'hc2b21bf7};
test_label[3722] = '{32'hc2b21bf7};
test_output[3722] = '{32'h432a42db};
/*############ DEBUG ############
test_input[29776:29783] = '{-98.7038536584, 62.6029462421, -57.4972072652, -28.9281000528, 81.2065402711, -4.47026247341, 4.31322932567, -89.0546172492};
test_label[3722] = '{-89.0546172492};
test_output[3722] = '{170.261157529};
############ END DEBUG ############*/
test_input[29784:29791] = '{32'hc23776df, 32'h41d0cf0b, 32'h4260e888, 32'hc1c854c7, 32'h4291ffc9, 32'hc2971b6e, 32'h42a2879f, 32'hbfd65659};
test_label[3723] = '{32'h42a2879f};
test_output[3723] = '{32'h3986e047};
/*############ DEBUG ############
test_input[29784:29791] = '{-45.86608687, 26.1010949494, 56.22708308, -25.041395157, 72.9995772158, -75.5535733408, 81.264888635, -1.67451014487};
test_label[3723] = '{81.264888635};
test_output[3723] = '{0.000257255707266};
############ END DEBUG ############*/
test_input[29792:29799] = '{32'hc25aec83, 32'h41854a70, 32'hc1b77f0c, 32'hc1c62aba, 32'hc1c64b1d, 32'hc294aae5, 32'h41bb2e9d, 32'h41bcbd03};
test_label[3724] = '{32'h41bcbd03};
test_output[3724] = '{32'h3f19e458};
/*############ DEBUG ############
test_input[29792:29799] = '{-54.7309682428, 16.6613458696, -22.9370340338, -24.7708619232, -24.7866769855, -74.3337767962, 23.3977609086, 23.5922915036};
test_label[3724] = '{23.5922915036};
test_output[3724] = '{0.601140475579};
############ END DEBUG ############*/
test_input[29800:29807] = '{32'h4234476f, 32'hc2a51501, 32'hc171b597, 32'hc2a425c5, 32'hbfb463e3, 32'hc293ecab, 32'hc06ca755, 32'h4264145c};
test_label[3725] = '{32'hc2a51501};
test_output[3725] = '{32'h430b8f98};
/*############ DEBUG ############
test_input[29800:29807] = '{45.0697611811, -82.5410226165, -15.106833106, -82.0737665775, -1.40929828934, -73.9622421149, -3.69771319909, 57.0198816908};
test_label[3725] = '{-82.5410226165};
test_output[3725] = '{139.560910766};
############ END DEBUG ############*/
test_input[29808:29815] = '{32'h42a9efe7, 32'hc2482938, 32'h41c0aaae, 32'h42c6f3f6, 32'hc22bb611, 32'h41c53052, 32'hc2c253e8, 32'hc28a5f8c};
test_label[3726] = '{32'hc2482938};
test_output[3726] = '{32'h43158449};
/*############ DEBUG ############
test_input[29808:29815] = '{84.9685563648, -50.0402531441, 24.0833395923, 99.4764825807, -42.9277989817, 24.6485930881, -97.1638818831, -69.1866168873};
test_label[3726] = '{-50.0402531441};
test_output[3726] = '{149.516736225};
############ END DEBUG ############*/
test_input[29816:29823] = '{32'hc1fb4e1b, 32'hc298305c, 32'hc1a8432b, 32'h41e79ba3, 32'h4285ce75, 32'h4233f342, 32'hc2acbf7c, 32'h427c40ce};
test_label[3727] = '{32'hc1a8432b};
test_output[3727] = '{32'h42afea24};
/*############ DEBUG ############
test_input[29816:29823] = '{-31.4131372735, -76.0944508123, -21.0327970066, 28.9509936346, 66.9032386144, 44.9875562308, -86.3739952371, 63.0632873397};
test_label[3727] = '{-21.0327970066};
test_output[3727] = '{87.9573025178};
############ END DEBUG ############*/
test_input[29824:29831] = '{32'hbf543baa, 32'hc20be7b5, 32'h42b508f4, 32'h4298c5cd, 32'hc1213e4a, 32'h428ee37c, 32'h4283c8c3, 32'h42162d5f};
test_label[3728] = '{32'h4298c5cd};
test_output[3728] = '{32'h4162193a};
/*############ DEBUG ############
test_input[29824:29831] = '{-0.829035406756, -34.9762748675, 90.5174859739, 76.3863278447, -10.0777077132, 71.444308493, 65.8921130022, 37.5443085102};
test_label[3728] = '{76.3863278447};
test_output[3728] = '{14.1311588638};
############ END DEBUG ############*/
test_input[29832:29839] = '{32'hc1e4eebc, 32'h415c6cd8, 32'h42c79e93, 32'hc20778da, 32'hbd25f672, 32'h42861357, 32'h3fdd082e, 32'h428d8281};
test_label[3729] = '{32'h415c6cd8};
test_output[3729] = '{32'h42ac10f8};
/*############ DEBUG ############
test_input[29832:29839] = '{-28.6165693718, 13.7765735039, 99.8097171176, -33.8680174323, -0.0405182316551, 67.0377701774, 1.72681217972, 70.754888125};
test_label[3729] = '{13.7765735039};
test_output[3729] = '{86.0331436137};
############ END DEBUG ############*/
test_input[29840:29847] = '{32'hc1885c47, 32'h421d3fd2, 32'h41b4d52c, 32'h4215ae24, 32'hc29097c4, 32'h42ae5e03, 32'hc2769155, 32'hc2a28b7e};
test_label[3730] = '{32'hc1885c47};
test_output[3730] = '{32'h42d07514};
/*############ DEBUG ############
test_input[29840:29847] = '{-17.0450576015, 39.3123244254, 22.604087463, 37.4200580856, -72.2964134684, 87.1836133299, -61.6419258438, -81.2724420086};
test_label[3730] = '{-17.0450576015};
test_output[3730] = '{104.228670931};
############ END DEBUG ############*/
test_input[29848:29855] = '{32'hc294b473, 32'h406deff7, 32'h425ffe5b, 32'hc23c926e, 32'h4188897f, 32'h422349ef, 32'hc2649716, 32'h4290b3e8};
test_label[3731] = '{32'h4188897f};
test_output[3731] = '{32'h425d2310};
/*############ DEBUG ############
test_input[29848:29855] = '{-74.3524435892, 3.71777137723, 55.998393666, -47.1429970942, 17.0671358458, 40.8222009986, -57.1475434112, 72.3513772138};
test_label[3731] = '{17.0671358458};
test_output[3731] = '{55.284241447};
############ END DEBUG ############*/
test_input[29856:29863] = '{32'h41382d6e, 32'hc183b90e, 32'hc2b8bdf7, 32'hc1bc09be, 32'hc0fd7cc8, 32'h42443330, 32'hc18d0181, 32'h42be2e9e};
test_label[3732] = '{32'h42be2e9e};
test_output[3732] = '{32'h80000000};
/*############ DEBUG ############
test_input[29856:29863] = '{11.5110908792, -16.4653592402, -92.371026373, -23.5047570235, -7.92148206407, 49.0499879996, -17.6257336661, 95.0910495606};
test_label[3732] = '{95.0910495606};
test_output[3732] = '{-0.0};
############ END DEBUG ############*/
test_input[29864:29871] = '{32'hc20f0973, 32'h42bd6152, 32'h422e5969, 32'h42975a33, 32'hc1918558, 32'hbf1bb34f, 32'h409d48cc, 32'h42bc976c};
test_label[3733] = '{32'h42975a33};
test_output[3733] = '{32'h419c3bcd};
/*############ DEBUG ############
test_input[29864:29871] = '{-35.7592285333, 94.6900797711, 43.5873158103, 75.6761739007, -18.1901086965, -0.608204793648, 4.91513631019, 94.2957465602};
test_label[3733] = '{75.6761739007};
test_output[3733] = '{19.5291991377};
############ END DEBUG ############*/
test_input[29872:29879] = '{32'hc2bda608, 32'h402025de, 32'h42530096, 32'h41e677ac, 32'hc2a0864f, 32'hc2972d49, 32'h42a84110, 32'hc2bcffdb};
test_label[3734] = '{32'h402025de};
test_output[3734] = '{32'h42a33fe1};
/*############ DEBUG ############
test_input[29872:29879] = '{-94.8242816548, 2.50231129546, 52.7505731337, 28.8084340379, -80.2623191609, -75.5884456974, 84.1270774092, -94.4997193271};
test_label[3734] = '{2.50231129546};
test_output[3734] = '{81.6247661138};
############ END DEBUG ############*/
test_input[29880:29887] = '{32'h41a34b77, 32'h428ea076, 32'hc1a8e6ca, 32'hc1e63f4c, 32'h4221434b, 32'hc2a063c5, 32'hc1d7cc55, 32'hc136edee};
test_label[3735] = '{32'h428ea076};
test_output[3735] = '{32'h291b8000};
/*############ DEBUG ############
test_input[29880:29887] = '{20.4118473774, 71.3134013494, -21.1126908757, -28.7809073186, 40.3157153813, -80.1948615664, -26.9747723654, -11.4330887252};
test_label[3735] = '{71.3134013494};
test_output[3735] = '{3.45279360658e-14};
############ END DEBUG ############*/
test_input[29888:29895] = '{32'hc2b4cb26, 32'hc1d6f843, 32'hc29670fd, 32'h41c756cd, 32'h42829cbb, 32'h3f317dc7, 32'h42250a3b, 32'h427eb2fd};
test_label[3736] = '{32'hc1d6f843};
test_output[3736] = '{32'h42b8b64b};
/*############ DEBUG ############
test_input[29888:29895] = '{-90.3967722032, -26.8712220463, -75.2206811156, 24.9173839359, 65.3061121487, 0.693325449099, 41.2599912721, 63.6747925807};
test_label[3736] = '{-26.8712220463};
test_output[3736] = '{92.3560418983};
############ END DEBUG ############*/
test_input[29896:29903] = '{32'hc2a3793c, 32'hc250a877, 32'hc255d0e6, 32'h420050d3, 32'h4191aa15, 32'h405b907b, 32'hc257dd68, 32'hc240ceb2};
test_label[3737] = '{32'h4191aa15};
test_output[3737] = '{32'h415def22};
/*############ DEBUG ############
test_input[29896:29903] = '{-81.7367877914, -52.1645181867, -53.45400342, 32.0789290268, 18.2080479485, 3.43069344551, -53.9662162432, -48.2018516858};
test_label[3737] = '{18.2080479485};
test_output[3737] = '{13.8708820244};
############ END DEBUG ############*/
test_input[29904:29911] = '{32'hc236fc63, 32'h4223a382, 32'h41fcd237, 32'hc1583d16, 32'hc1f45527, 32'h422422ac, 32'hc16350c7, 32'hc2b099ca};
test_label[3738] = '{32'h4223a382};
test_output[3738] = '{32'h3f41d860};
/*############ DEBUG ############
test_input[29904:29911] = '{-45.7464714693, 40.9096765228, 31.602643989, -13.5149140113, -30.5415783451, 41.033859812, -14.2072209724, -88.3003724093};
test_label[3738] = '{40.9096765228};
test_output[3738] = '{0.757207849949};
############ END DEBUG ############*/
test_input[29912:29919] = '{32'h422a10d8, 32'h42944464, 32'h4150ec9b, 32'h423cfa03, 32'h426b0c34, 32'hc2240e58, 32'h42bb8aba, 32'hc228a2c8};
test_label[3739] = '{32'h42944464};
test_output[3739] = '{32'h419d1959};
/*############ DEBUG ############
test_input[29912:29919] = '{42.5164496589, 74.1335716649, 13.0577650706, 47.2441510506, 58.7619179981, -41.0140072031, 93.7709475533, -42.1589679323};
test_label[3739] = '{74.1335716649};
test_output[3739] = '{19.6373758913};
############ END DEBUG ############*/
test_input[29920:29927] = '{32'h42ad43a1, 32'h41b5a8db, 32'hc24f2a84, 32'h40e84066, 32'hc183a1e8, 32'h40c8f35c, 32'h42b6e5c3, 32'hc2bdd63a};
test_label[3740] = '{32'h41b5a8db};
test_output[3740] = '{32'h42897fad};
/*############ DEBUG ############
test_input[29920:29927] = '{86.632090628, 22.7074488568, -51.7915183643, 7.25786135988, -16.4540560113, 6.27970683283, 91.4487525658, -94.9184091019};
test_label[3740] = '{22.7074488568};
test_output[3740] = '{68.7493648898};
############ END DEBUG ############*/
test_input[29928:29935] = '{32'hc2948f14, 32'hc2b30a52, 32'hc27c94ec, 32'hc287247b, 32'h41d59c42, 32'hc2823d69, 32'h42ad1168, 32'hc2703c94};
test_label[3741] = '{32'hc2948f14};
test_output[3741] = '{32'h4320d03e};
/*############ DEBUG ############
test_input[29928:29935] = '{-74.2794505187, -89.5201593782, -63.1454324371, -67.5712538486, 26.7012982963, -65.1199418126, 86.5339931353, -60.059156666};
test_label[3741] = '{-74.2794505187};
test_output[3741] = '{160.813443654};
############ END DEBUG ############*/
test_input[29936:29943] = '{32'hc28e66cf, 32'h428f839f, 32'h428ef3df, 32'h42961cee, 32'h42490054, 32'h41ebc160, 32'h428c80a9, 32'h4134afce};
test_label[3742] = '{32'h428f839f};
test_output[3742] = '{32'h4057abb3};
/*############ DEBUG ############
test_input[29936:29943] = '{-71.2007969502, 71.7570745622, 71.4763137828, 75.0565068276, 50.2503190529, 29.4694215039, 70.2512875474, 11.2929206339};
test_label[3742] = '{71.7570745622};
test_output[3742] = '{3.36985469517};
############ END DEBUG ############*/
test_input[29944:29951] = '{32'hc23545c9, 32'h42c0875f, 32'h4254138a, 32'hc25e716d, 32'hc2016cc5, 32'h428a2180, 32'h42c5965a, 32'hc2788479};
test_label[3743] = '{32'hc23545c9};
test_output[3743] = '{32'h43103042};
/*############ DEBUG ############
test_input[29944:29951] = '{-45.3181478667, 96.2643998181, 53.0190804627, -55.610768225, -32.3562200518, 69.0654268817, 98.7936559545, -62.1293670135};
test_label[3743] = '{-45.3181478667};
test_output[3743] = '{144.188503993};
############ END DEBUG ############*/
test_input[29952:29959] = '{32'hc207d2e6, 32'hc119f800, 32'hc221a241, 32'h42b7190e, 32'h41c65779, 32'hc19ba60c, 32'hc2911b59, 32'hc18708b8};
test_label[3744] = '{32'hc19ba60c};
test_output[3744] = '{32'h42de0291};
/*############ DEBUG ############
test_input[29952:29959] = '{-33.9559542308, -9.62304695593, -40.4084495431, 91.5489323472, 24.7927107453, -19.4560776682, -72.5534156725, -16.8792570053};
test_label[3744] = '{-19.4560776682};
test_output[3744] = '{111.005010015};
############ END DEBUG ############*/
test_input[29960:29967] = '{32'hc1cd9674, 32'h428e1eff, 32'hc08260cc, 32'h42c3568f, 32'h42878f19, 32'h41e2e129, 32'hc2a33a3c, 32'hc26ac6c4};
test_label[3745] = '{32'h428e1eff};
test_output[3745] = '{32'h41d4de3f};
/*############ DEBUG ############
test_input[29960:29967] = '{-25.6984636487, 71.0605410038, -4.07431596569, 97.6690600475, 67.7794888381, 28.3599412101, -81.6137422193, -58.6941064283};
test_label[3745] = '{71.0605410038};
test_output[3745] = '{26.6085190437};
############ END DEBUG ############*/
test_input[29968:29975] = '{32'h424f65b6, 32'h3fed1650, 32'h42a73e00, 32'h423ad9cf, 32'hc294a3e2, 32'h42093f3c, 32'hc2212b8f, 32'hc1d9817a};
test_label[3746] = '{32'h42093f3c};
test_output[3746] = '{32'h42453cc5};
/*############ DEBUG ############
test_input[29968:29975] = '{51.849327807, 1.85224346447, 83.6210941534, 46.7127032068, -74.3200869396, 34.311750479, -40.2925393186, -27.1882213442};
test_label[3746] = '{34.311750479};
test_output[3746] = '{49.3093436745};
############ END DEBUG ############*/
test_input[29976:29983] = '{32'h42982aa7, 32'h426c1ff1, 32'h42b8c7ca, 32'hc29f908a, 32'h4056e1f8, 32'h42709c69, 32'hc1201147, 32'hc1803212};
test_label[3747] = '{32'h42982aa7};
test_output[3747] = '{32'h4182748c};
/*############ DEBUG ############
test_input[29976:29983] = '{76.0833089983, 59.0311910914, 92.3902160804, -79.782301197, 3.35754199846, 60.1527443377, -10.0042183258, -16.0244492505};
test_label[3747] = '{76.0833089983};
test_output[3747] = '{16.3069071648};
############ END DEBUG ############*/
test_input[29984:29991] = '{32'h41dea100, 32'hc1b516ab, 32'h417797f0, 32'hc1cbe306, 32'hc279632b, 32'hc094c009, 32'h4279c4b2, 32'h42b0cf74};
test_label[3748] = '{32'h417797f0};
test_output[3748] = '{32'h4291dc76};
/*############ DEBUG ############
test_input[29984:29991] = '{27.8286134316, -22.6360687032, 15.4745941797, -25.4858515129, -62.3468434797, -4.64844197642, 62.4420837476, 88.4051798746};
test_label[3748] = '{15.4745941797};
test_output[3748] = '{72.9305856949};
############ END DEBUG ############*/
test_input[29992:29999] = '{32'hc27863d2, 32'h41fc5396, 32'hc0cdec37, 32'hc2ab4d96, 32'hc2b6739c, 32'h42ac3031, 32'h427e4ab8, 32'hc2428d1c};
test_label[3749] = '{32'h427e4ab8};
test_output[3749] = '{32'h41b42b56};
/*############ DEBUG ############
test_input[29992:29999] = '{-62.0974812614, 31.5408136587, -6.43508463301, -85.6515316046, -91.2257965555, 86.0941274015, 63.5729678887, -48.6378005647};
test_label[3749] = '{63.5729678887};
test_output[3749] = '{22.521159513};
############ END DEBUG ############*/
test_input[30000:30007] = '{32'h419af085, 32'h4292b9d2, 32'h421cdeb5, 32'hc2a4d7d4, 32'h42884d77, 32'hc2492caa, 32'hc03b51b9, 32'hc29d4d66};
test_label[3750] = '{32'hc2492caa};
test_output[3750] = '{32'h42f752f0};
/*############ DEBUG ############
test_input[30000:30007] = '{19.367441506, 73.3629279102, 39.2174869864, -82.4215393535, 68.1512974262, -50.2936185106, -2.92686307255, -78.6511665404};
test_label[3750] = '{-50.2936185106};
test_output[3750] = '{123.661984384};
############ END DEBUG ############*/
test_input[30008:30015] = '{32'hc2ba3d02, 32'hc2727ba8, 32'h42590b29, 32'h423d2a47, 32'hc102af62, 32'h40fa86fd, 32'h42c39a5c, 32'hc29cf8cd};
test_label[3751] = '{32'h42590b29};
test_output[3751] = '{32'h422e298f};
/*############ DEBUG ############
test_input[30008:30015] = '{-93.11915466, -60.6207591241, 54.2608995968, 47.2912874069, -8.16781824413, 7.82897829657, 97.8014842273, -78.4859412982};
test_label[3751] = '{54.2608995968};
test_output[3751] = '{43.5405846305};
############ END DEBUG ############*/
test_input[30016:30023] = '{32'h4281128f, 32'h411ff66f, 32'h42a922ab, 32'h42bc0d0a, 32'hc2b1c507, 32'hc2a98acb, 32'h4251ad55, 32'h42c78b56};
test_label[3752] = '{32'h42c78b56};
test_output[3752] = '{32'h3b50f718};
/*############ DEBUG ############
test_input[30016:30023] = '{64.5362437255, 9.99766424598, 84.5677108815, 94.0254698171, -88.884821631, -84.7710835084, 52.419270779, 99.7721403331};
test_label[3752] = '{99.7721403331};
test_output[3752] = '{0.00318855596794};
############ END DEBUG ############*/
test_input[30024:30031] = '{32'h4235164c, 32'hbf45dde1, 32'h425da0c9, 32'h41f4e9ff, 32'hc1afb85c, 32'hc1e899a1, 32'hc2834714, 32'h4280129d};
test_label[3753] = '{32'h4235164c};
test_output[3753] = '{32'h41961e39};
/*############ DEBUG ############
test_input[30024:30031] = '{45.2717737032, -0.772916846983, 55.4070155165, 30.614255963, -21.9650188111, -29.0750131841, -65.6388240782, 64.0363522056};
test_label[3753] = '{45.2717737032};
test_output[3753] = '{18.7647572767};
############ END DEBUG ############*/
test_input[30032:30039] = '{32'h42b45221, 32'h42c79ae8, 32'hc28cd210, 32'h41d23ebd, 32'hc239de35, 32'h42907b70, 32'hc294a882, 32'hc198b858};
test_label[3754] = '{32'h42b45221};
test_output[3754] = '{32'h411a4678};
/*############ DEBUG ############
test_input[30032:30039] = '{90.1604109371, 99.8025506252, -70.4102811274, 26.2806342203, -46.4670008298, 72.2410888497, -74.3291190365, -19.0900110568};
test_label[3754] = '{90.1604109371};
test_output[3754] = '{9.64220461993};
############ END DEBUG ############*/
test_input[30040:30047] = '{32'hc2b11620, 32'h427122a2, 32'hc24a4687, 32'h4208df67, 32'hc20a800e, 32'hc124769f, 32'hc14b6263, 32'hc2127e42};
test_label[3755] = '{32'hc2127e42};
test_output[3755] = '{32'h42c1d072};
/*############ DEBUG ############
test_input[30040:30047] = '{-88.5432139848, 60.2838200832, -50.5688753624, 34.2181647632, -34.6250540981, -10.2789603072, -12.711520089, -36.623298332};
test_label[3755] = '{-36.623298332};
test_output[3755] = '{96.9071184152};
############ END DEBUG ############*/
test_input[30048:30055] = '{32'hc27bffde, 32'hc1c4a349, 32'h42c29879, 32'hc29254d9, 32'hc1d48614, 32'hc2a734c9, 32'hc289a907, 32'hc01d2861};
test_label[3756] = '{32'hc1d48614};
test_output[3756] = '{32'h42f7b9fe};
/*############ DEBUG ############
test_input[30048:30055] = '{-62.9998721607, -24.5797292341, 97.2977950562, -73.1657218346, -26.5654681306, -83.6030957616, -68.8301318887, -2.45558954976};
test_label[3756] = '{-26.5654681306};
test_output[3756] = '{123.863263187};
############ END DEBUG ############*/
test_input[30056:30063] = '{32'hc254ae53, 32'h41c25e21, 32'h429fc187, 32'hc2700cdc, 32'hc16944d9, 32'hc2057d73, 32'h42a25202, 32'hc29ef601};
test_label[3757] = '{32'h41c25e21};
test_output[3757] = '{32'h42646fad};
/*############ DEBUG ############
test_input[30056:30063] = '{-53.1702373467, 24.2959615883, 79.8779793634, -60.0125589015, -14.5793082558, -33.3725097424, 81.1601698876, -79.4804753152};
test_label[3757] = '{24.2959615883};
test_output[3757] = '{57.1090577006};
############ END DEBUG ############*/
test_input[30064:30071] = '{32'h4186cec9, 32'h4180b87a, 32'h415e9e2f, 32'h429719b8, 32'h42c6bbd3, 32'h42a31e1b, 32'h40a92b84, 32'h4299ed71};
test_label[3758] = '{32'h4186cec9};
test_output[3758] = '{32'h42a50821};
/*############ DEBUG ############
test_input[30064:30071] = '{16.8509694259, 16.0900767612, 13.9136188706, 75.5502284557, 99.3668469833, 81.5587960547, 5.2865620914, 76.9637528376};
test_label[3758] = '{16.8509694259};
test_output[3758] = '{82.5158775761};
############ END DEBUG ############*/
test_input[30072:30079] = '{32'hc25bb953, 32'hc1073db4, 32'h428a9a78, 32'h4227090b, 32'hc1ae933b, 32'hc26ac031, 32'h412b449f, 32'hc146ab70};
test_label[3759] = '{32'hc26ac031};
test_output[3759] = '{32'h42fffa90};
/*############ DEBUG ############
test_input[30072:30079] = '{-54.9309810256, -8.45256420875, 69.3016962533, 41.7588324348, -21.8218891563, -58.6876865395, 10.7042533173, -12.4168552053};
test_label[3759] = '{-58.6876865395};
test_output[3759] = '{127.989382793};
############ END DEBUG ############*/
test_input[30080:30087] = '{32'h429a82b2, 32'h42600407, 32'hc2418b6f, 32'hc28ec3c2, 32'h42898040, 32'h4251c489, 32'h41badcb8, 32'h42647859};
test_label[3760] = '{32'h4251c489};
test_output[3760] = '{32'h41c68221};
/*############ DEBUG ############
test_input[30080:30087] = '{77.2552647924, 56.003934582, -48.386165444, -71.3823425456, 68.75048997, 52.4419276641, 23.3577723071, 57.1175263041};
test_label[3760] = '{52.4419276641};
test_output[3760] = '{24.8135396094};
############ END DEBUG ############*/
test_input[30088:30095] = '{32'h42015999, 32'hc294206f, 32'hc16397ab, 32'h4225f525, 32'hc238a8dc, 32'h3fe4622c, 32'h427e2ad1, 32'hc1c94896};
test_label[3761] = '{32'h4225f525};
test_output[3761] = '{32'h41b06b58};
/*############ DEBUG ############
test_input[30088:30095] = '{32.3374993365, -74.0633493937, -14.2245286576, 41.4893974439, -46.1649007208, 1.78424592689, 63.5418113759, -25.1604422964};
test_label[3761] = '{41.4893974439};
test_output[3761] = '{22.0524139322};
############ END DEBUG ############*/
test_input[30096:30103] = '{32'hc293191e, 32'h429e96a2, 32'h42173c87, 32'hc25fe525, 32'hc22e71f1, 32'hc20688e7, 32'hc28549c9, 32'h42b26c8a};
test_label[3762] = '{32'hc20688e7};
test_output[3762] = '{32'h42f5b104};
/*############ DEBUG ############
test_input[30096:30103] = '{-73.5490566751, 79.2942019413, 37.8091082277, -55.973773539, -43.6112725022, -33.6336947671, -66.6441095293, 89.2119917096};
test_label[3762] = '{-33.6336947671};
test_output[3762] = '{122.845735765};
############ END DEBUG ############*/
test_input[30104:30111] = '{32'h42977647, 32'hc1e4a0bd, 32'h4075268f, 32'h42187123, 32'hc2c0f994, 32'hc28772f3, 32'hc2a41035, 32'hc2a57766};
test_label[3763] = '{32'h4075268f};
test_output[3763] = '{32'h428fcd13};
/*############ DEBUG ############
test_input[30104:30111] = '{75.7310138462, -28.5784863229, 3.83047842351, 38.1104843486, -96.4874581379, -67.7245075091, -82.0316535122, -82.7332018121};
test_label[3763] = '{3.83047842351};
test_output[3763] = '{71.9005354227};
############ END DEBUG ############*/
test_input[30112:30119] = '{32'hc2937771, 32'h428b168e, 32'h42b27834, 32'hc02d95f9, 32'hc1fa4a16, 32'h41df6231, 32'h427da27c, 32'hc2956bf1};
test_label[3764] = '{32'h42b27834};
test_output[3764] = '{32'h314165b5};
/*############ DEBUG ############
test_input[30112:30119] = '{-73.7332830455, 69.5440538187, 89.2347683124, -2.7122786009, -31.286174682, 27.9229447828, 63.4086772488, -74.7108206079};
test_label[3764] = '{89.2347683124};
test_output[3764] = '{2.81430090739e-09};
############ END DEBUG ############*/
test_input[30120:30127] = '{32'h41e659bd, 32'h4227be05, 32'h3f696a14, 32'h42922fc0, 32'h42c178e9, 32'hc2996c23, 32'h42a520ef, 32'h41629c39};
test_label[3765] = '{32'hc2996c23};
test_output[3765] = '{32'h432d7286};
/*############ DEBUG ############
test_input[30120:30127] = '{28.7938167317, 41.9355649392, 0.91177489993, 73.0932605407, 96.7361495207, -76.7112029243, 82.5643221211, 14.1631405514};
test_label[3765] = '{-76.7112029243};
test_output[3765] = '{173.447353145};
############ END DEBUG ############*/
test_input[30128:30135] = '{32'h423280e8, 32'h41d9ffbb, 32'hc22d75fb, 32'hbf067bae, 32'h42887199, 32'h41cd62f4, 32'h421bd158, 32'h429bbc26};
test_label[3766] = '{32'h423280e8};
test_output[3766] = '{32'h4204f775};
/*############ DEBUG ############
test_input[30128:30135] = '{44.62588657, 27.2498691916, -43.3652162524, -0.525324715795, 68.2218678416, 25.6733164395, 38.954438242, 77.8674796559};
test_label[3766] = '{44.62588657};
test_output[3766] = '{33.2416577927};
############ END DEBUG ############*/
test_input[30136:30143] = '{32'h4178b261, 32'h425dedce, 32'h41f761a1, 32'h41a35296, 32'hc230581c, 32'h404f0cb6, 32'h421f4131, 32'hc1d5c039};
test_label[3767] = '{32'h425dedce};
test_output[3767] = '{32'h342856ef};
/*############ DEBUG ############
test_input[30136:30143] = '{15.5435491379, 55.4822327944, 30.922669692, 20.4153256039, -44.0860450524, 3.23515070768, 39.8136631434, -26.7188586697};
test_label[3767] = '{55.4822327944};
test_output[3767] = '{1.56778459736e-07};
############ END DEBUG ############*/
test_input[30144:30151] = '{32'h4252cb02, 32'h4264b4bd, 32'hc1b7666b, 32'h424fa545, 32'hc29fd1c6, 32'h4258e5f9, 32'h4231af8e, 32'h42a09e49};
test_label[3768] = '{32'h4258e5f9};
test_output[3768] = '{32'h41d0ad32};
/*############ DEBUG ############
test_input[30144:30151] = '{52.6982510798, 57.176500957, -22.9250084218, 51.9113952293, -79.9097111443, 54.2245825312, 44.4214386338, 80.3091498783};
test_label[3768] = '{54.2245825312};
test_output[3768] = '{26.0845673472};
############ END DEBUG ############*/
test_input[30152:30159] = '{32'h411f29dd, 32'h42a3efd6, 32'hc2a007cd, 32'h4195a977, 32'h4288614e, 32'h41e79af8, 32'hc20c9672, 32'h423b5e0c};
test_label[3769] = '{32'hc20c9672};
test_output[3769] = '{32'h42ea3b0f};
/*############ DEBUG ############
test_input[30152:30159] = '{9.94772005778, 81.9684292836, -80.0152348811, 18.7077473858, 68.190045861, 28.9506686686, -35.1469200573, 46.8418419836};
test_label[3769] = '{-35.1469200573};
test_output[3769] = '{117.115350379};
############ END DEBUG ############*/
test_input[30160:30167] = '{32'hc2b46723, 32'h42ad2062, 32'hc226a8a7, 32'hc290ab6b, 32'hc2858e48, 32'hc0fc82c2, 32'hc246bcf1, 32'hc2a0f647};
test_label[3770] = '{32'hc246bcf1};
test_output[3770] = '{32'h43083f6d};
/*############ DEBUG ############
test_input[30160:30167] = '{-90.2014372479, 86.5632463904, -41.6646996339, -72.334798483, -66.7778934735, -7.89096162143, -49.6845112822, -80.4810075279};
test_label[3770] = '{-49.6845112822};
test_output[3770] = '{136.247757673};
############ END DEBUG ############*/
test_input[30168:30175] = '{32'hc2b56483, 32'h42524d0f, 32'h429b1d17, 32'hc270e539, 32'h42986aeb, 32'hc19f396e, 32'hc229f18d, 32'hc217d7ce};
test_label[3771] = '{32'hc270e539};
test_output[3771] = '{32'h430a02f7};
/*############ DEBUG ############
test_input[30168:30175] = '{-90.6963150102, 52.5752520337, 77.5568174218, -60.2238487634, 76.2088260878, -19.9030421261, -42.4858904403, -37.9607469065};
test_label[3771] = '{-60.2238487634};
test_output[3771] = '{138.011588611};
############ END DEBUG ############*/
test_input[30176:30183] = '{32'h42900400, 32'h42a9e175, 32'hc10e6f1e, 32'hc225bf60, 32'hc2b935e6, 32'h42c1b113, 32'hc235624c, 32'h418ac723};
test_label[3772] = '{32'h42c1b113};
test_output[3772] = '{32'h36e29941};
/*############ DEBUG ############
test_input[30176:30183] = '{72.0078134531, 84.9403464937, -8.90212817271, -41.4368910094, -92.6052691371, 96.8458446545, -45.3459917335, 17.347233986};
test_label[3772] = '{96.8458446545};
test_output[3772] = '{6.75316604585e-06};
############ END DEBUG ############*/
test_input[30184:30191] = '{32'hc0be8204, 32'h42c19e22, 32'hc28d4eb7, 32'h41efe8c1, 32'hc1d66dce, 32'hc25e195d, 32'h42770a24, 32'hc2a1cbcf};
test_label[3773] = '{32'h42770a24};
test_output[3773] = '{32'h420c3220};
/*############ DEBUG ############
test_input[30184:30191] = '{-5.95337101725, 96.8088545567, -70.6537370748, 29.9886495529, -26.8036157813, -55.5247696577, 61.7599044597, -80.8980614033};
test_label[3773] = '{61.7599044597};
test_output[3773] = '{35.048950097};
############ END DEBUG ############*/
test_input[30192:30199] = '{32'hc261b00f, 32'hc16f6c92, 32'hc2a9c634, 32'hc28381fc, 32'h42c54c18, 32'hc272053a, 32'hc255691e, 32'h42c2ec26};
test_label[3774] = '{32'hc261b00f};
test_output[3774] = '{32'h431b5637};
/*############ DEBUG ############
test_input[30192:30199] = '{-56.4219338586, -14.9640068674, -84.8871160752, -65.7538771933, 98.6486242629, -60.5051057634, -53.3526542905, 97.4612291543};
test_label[3774] = '{-56.4219338586};
test_output[3774] = '{155.336772473};
############ END DEBUG ############*/
test_input[30200:30207] = '{32'h42ab5e3d, 32'h41c2075f, 32'h428f085a, 32'h42ad0422, 32'h42693ac0, 32'h3f7b443a, 32'h4253afe7, 32'hc2289317};
test_label[3775] = '{32'h42ab5e3d};
test_output[3775] = '{32'h3f980787};
/*############ DEBUG ############
test_input[30200:30207] = '{85.6840627009, 24.2535989671, 71.5163144978, 86.5080742526, 58.3073743105, 0.981509786472, 52.9217811403, -42.1436418419};
test_label[3775] = '{85.6840627009};
test_output[3775] = '{1.18772971522};
############ END DEBUG ############*/
test_input[30208:30215] = '{32'h418d81e1, 32'h42c74db6, 32'h3e4b8b02, 32'hc293f232, 32'hc2872460, 32'h41393b42, 32'h42c3b9ba, 32'h3ecdb1da};
test_label[3776] = '{32'h41393b42};
test_output[3776] = '{32'h42b0756e};
/*############ DEBUG ############
test_input[30208:30215] = '{17.6884166264, 99.6517818511, 0.198772464988, -73.9730356114, -67.5710437474, 11.5769671255, 97.8627469692, 0.401747539014};
test_label[3776] = '{11.5769671255};
test_output[3776] = '{88.229355087};
############ END DEBUG ############*/
test_input[30216:30223] = '{32'hc20ffd0c, 32'hc28f579f, 32'hc29366c0, 32'hc123e8f4, 32'h42764729, 32'hc112f8c7, 32'hc121f063, 32'h429322ff};
test_label[3777] = '{32'hc121f063};
test_output[3777] = '{32'h42a7610c};
/*############ DEBUG ############
test_input[30216:30223] = '{-35.9971146418, -71.6711374618, -73.7006813425, -10.244372904, 61.5694927918, -9.18573705079, -10.1211886146, 73.5683509628};
test_label[3777] = '{-10.1211886146};
test_output[3777] = '{83.6895457286};
############ END DEBUG ############*/
test_input[30224:30231] = '{32'h42275d82, 32'h4269bf8d, 32'hbfdc84c5, 32'h40c95333, 32'hc23a9760, 32'h42094f66, 32'h425da6bd, 32'hc2a987e0};
test_label[3778] = '{32'hbfdc84c5};
test_output[3778] = '{32'h4270d44a};
/*############ DEBUG ############
test_input[30224:30231] = '{41.8413168914, 58.4370613561, -1.72280183734, 6.29140626604, -46.6478276217, 34.3275357841, 55.4128319244, -84.7653810393};
test_label[3778] = '{-1.72280183734};
test_output[3778] = '{60.2073146666};
############ END DEBUG ############*/
test_input[30232:30239] = '{32'hc178be07, 32'hc151f11b, 32'hc26c3e97, 32'hc23cf2b9, 32'h42b12222, 32'h40e1e0ae, 32'h41612edd, 32'h4104fb7d};
test_label[3779] = '{32'h41612edd};
test_output[3779] = '{32'h4294fc47};
/*############ DEBUG ############
test_input[30232:30239] = '{-15.5463930344, -13.1213638502, -59.0611232689, -47.237033449, 88.5666693349, 7.05867659918, 14.0739409649, 8.31139809111};
test_label[3779] = '{14.0739409649};
test_output[3779] = '{74.49272837};
############ END DEBUG ############*/
test_input[30240:30247] = '{32'h425d61fc, 32'h4192c162, 32'hc290772b, 32'hc1996e08, 32'hc21e75d8, 32'h42a2ec1b, 32'h4279f03b, 32'hc1dd2328};
test_label[3780] = '{32'h42a2ec1b};
test_output[3780] = '{32'h31c53c7b};
/*############ DEBUG ############
test_input[30240:30247] = '{55.3456873771, 18.3444254735, -72.2327502363, -19.1787267035, -39.6150802581, 81.4611408543, 62.4845984867, -27.6421662408};
test_label[3780] = '{81.4611408543};
test_output[3780] = '{5.74033044969e-09};
############ END DEBUG ############*/
test_input[30248:30255] = '{32'hc0cd9b42, 32'h429811dd, 32'h40bf516f, 32'hc2795d33, 32'hc28343d4, 32'hc2023396, 32'hc1aabd1d, 32'h414fde6d};
test_label[3781] = '{32'hc2795d33};
test_output[3781] = '{32'h430a603b};
/*############ DEBUG ############
test_input[30248:30255] = '{-6.42520250627, 76.03489243, 5.97869052297, -62.3410137323, -65.6324741559, -32.5503780568, -21.342340482, 12.991802715};
test_label[3781] = '{-62.3410137323};
test_output[3781] = '{138.375906162};
############ END DEBUG ############*/
test_input[30256:30263] = '{32'hc1a1fbf8, 32'hc247605f, 32'hc2aa7ccd, 32'h421f40db, 32'hc16c47ef, 32'h428e15aa, 32'h41c5f85d, 32'hbedbca4a};
test_label[3782] = '{32'hbedbca4a};
test_output[3782] = '{32'h428ef174};
/*############ DEBUG ############
test_input[30256:30263] = '{-20.2480324857, -49.844112713, -85.2437543727, 39.8133369756, -14.7675617662, 71.0423088835, 24.7462711923, -0.429277713979};
test_label[3782] = '{-0.429277713979};
test_output[3782] = '{71.4715865975};
############ END DEBUG ############*/
test_input[30264:30271] = '{32'hc297f80b, 32'hc2c74894, 32'h426dea5d, 32'hc1f4058b, 32'h41f0f26e, 32'hc28ba64d, 32'hc1d546fc, 32'h42bb780f};
test_label[3783] = '{32'h41f0f26e};
test_output[3783] = '{32'h427e76e7};
/*############ DEBUG ############
test_input[30264:30271] = '{-75.9844622809, -99.6417569053, 59.4788706258, -30.5027071862, 30.1183742442, -69.8248039187, -26.6596599719, 93.7344888395};
test_label[3783] = '{30.1183742442};
test_output[3783] = '{63.6161145952};
############ END DEBUG ############*/
test_input[30272:30279] = '{32'h42a378f7, 32'h42201c0d, 32'hc1506a8c, 32'hc20c0324, 32'hbf9ddc60, 32'h421ba3cf, 32'hc1b650d9, 32'h4281ea79};
test_label[3784] = '{32'hc1b650d9};
test_output[3784] = '{32'h42d10d2d};
/*############ DEBUG ############
test_input[30272:30279] = '{81.7362568475, 40.0273947132, -13.0260123747, -35.0030688259, -1.23328779888, 38.9099690064, -22.7894756024, 64.9579557151};
test_label[3784] = '{-22.7894756024};
test_output[3784] = '{104.525732502};
############ END DEBUG ############*/
test_input[30280:30287] = '{32'hc159db22, 32'hc12b5af9, 32'h4224ba40, 32'h42ab264c, 32'hc210bb82, 32'h413edc0c, 32'hc0b22126, 32'h423ba9f1};
test_label[3785] = '{32'hc12b5af9};
test_output[3785] = '{32'h42c091ac};
/*############ DEBUG ############
test_input[30280:30287] = '{-13.6159992343, -10.7097104078, 41.1818848947, 85.5748021316, -36.1831141573, 11.9287224071, -5.56654644606, 46.9159583001};
test_label[3785] = '{-10.7097104078};
test_output[3785] = '{96.2845125394};
############ END DEBUG ############*/
test_input[30288:30295] = '{32'h42250cf4, 32'hc143ffa4, 32'hc2114428, 32'hc1f57908, 32'hc130d8ea, 32'hc2bcc1ea, 32'hc121b419, 32'hc293ff23};
test_label[3786] = '{32'hc2bcc1ea};
test_output[3786] = '{32'h4307a432};
/*############ DEBUG ############
test_input[30288:30295] = '{41.2626502614, -12.2499124859, -36.3165595517, -30.6840981502, -11.0529574, -94.3787355355, -10.1064690854, -73.9983133408};
test_label[3786] = '{-94.3787355355};
test_output[3786] = '{135.641385797};
############ END DEBUG ############*/
test_input[30296:30303] = '{32'hc28d94dc, 32'hc29120a1, 32'h41f7548c, 32'hc258c07d, 32'hc284c3b7, 32'h4287e0c8, 32'h4241588e, 32'h417cd4b3};
test_label[3787] = '{32'h4287e0c8};
test_output[3787] = '{32'h3152c436};
/*############ DEBUG ############
test_input[30296:30303] = '{-70.7907386642, -72.5637305924, 30.9162832005, -54.1879769708, -66.3822568037, 67.9390270373, 48.3364791594, 15.8019282014};
test_label[3787] = '{67.9390270373};
test_output[3787] = '{3.06705550317e-09};
############ END DEBUG ############*/
test_input[30304:30311] = '{32'hc1bb553d, 32'h4215c923, 32'h4140a9aa, 32'h4284725f, 32'h423caa51, 32'h423406a6, 32'h41960a2d, 32'hc2aaa4c3};
test_label[3788] = '{32'h41960a2d};
test_output[3788] = '{32'h423ddfa7};
/*############ DEBUG ############
test_input[30304:30311] = '{-23.4166194749, 37.4464243089, 12.0414223591, 66.2233781616, 47.1663233321, 45.0064926113, 18.7549677123, -85.3218020317};
test_label[3788] = '{18.7549677123};
test_output[3788] = '{47.4684104552};
############ END DEBUG ############*/
test_input[30312:30319] = '{32'h42a06b5d, 32'hc21e6657, 32'hc23976f6, 32'hc21eb38a, 32'hc280b68f, 32'h429a7fd8, 32'h4284b0e0, 32'hc25705cc};
test_label[3789] = '{32'hc23976f6};
test_output[3789] = '{32'h42fd40b6};
/*############ DEBUG ############
test_input[30312:30319] = '{80.2096943461, -39.5999407736, -46.3661722156, -39.675332304, -64.3565628633, 77.2496961073, 66.3454569064, -53.7556608217};
test_label[3789] = '{-46.3661722156};
test_output[3789] = '{126.626388522};
############ END DEBUG ############*/
test_input[30320:30327] = '{32'h4266b928, 32'hc2abeb6f, 32'h42b7c0a9, 32'h41b9aa17, 32'hc2872728, 32'hc297bf7f, 32'hc22bbad9, 32'h42a6595d};
test_label[3790] = '{32'h41b9aa17};
test_output[3790] = '{32'h42895639};
/*############ DEBUG ############
test_input[30320:30327] = '{57.6808149767, -85.9598350332, 91.87628659, 23.2080516295, -67.576474864, -75.8740164031, -42.9324667399, 83.1745402193};
test_label[3790] = '{23.2080516295};
test_output[3790] = '{68.6684012418};
############ END DEBUG ############*/
test_input[30328:30335] = '{32'hc2c4819d, 32'hc2846515, 32'hc20c928a, 32'h42aeecf5, 32'hc2bbe8aa, 32'h42bf76b4, 32'hc1568726, 32'h423948fb};
test_label[3791] = '{32'hc2c4819d};
test_output[3791] = '{32'h4341fc39};
/*############ DEBUG ############
test_input[30328:30335] = '{-98.2531483617, -66.1974259464, -35.1431034675, 87.4628071396, -93.9544186416, 95.7318386108, -13.4079948045, 46.3212701451};
test_label[3791] = '{-98.2531483617};
test_output[3791] = '{193.985243273};
############ END DEBUG ############*/
test_input[30336:30343] = '{32'h42893aab, 32'h42b0a6ca, 32'hc1e27021, 32'h41addbcb, 32'h42c067d0, 32'h428cdc4e, 32'h41869059, 32'hc2a163fc};
test_label[3792] = '{32'h41869059};
test_output[3792] = '{32'h429ec3ec};
/*############ DEBUG ############
test_input[30336:30343] = '{68.6145890477, 88.3257633029, -28.3047506897, 21.7323206052, 96.2027615084, 70.4302826949, 16.8204818972, -80.6952801774};
test_label[3792] = '{16.8204818972};
test_output[3792] = '{79.3826589094};
############ END DEBUG ############*/
test_input[30344:30351] = '{32'h40e84512, 32'hc27bda71, 32'h426d5ac7, 32'h40f93616, 32'h426cff3f, 32'hc05ca7f4, 32'hc22b479b, 32'hc2a5f78e};
test_label[3793] = '{32'h40f93616};
test_output[3793] = '{32'h4250cd0e};
/*############ DEBUG ############
test_input[30344:30351] = '{7.25843139611, -62.9633210364, 59.3386492931, 7.78785220859, 59.2492643185, -3.44775112794, -42.8199271574, -82.9835055874};
test_label[3793] = '{7.78785220859};
test_output[3793] = '{52.2002501547};
############ END DEBUG ############*/
test_input[30352:30359] = '{32'h42b2a0a2, 32'hc1e8bcee, 32'hc18d122e, 32'hc2710bac, 32'h4134abb2, 32'h42b7fd92, 32'hc18580e2, 32'hc2a14ef9};
test_label[3794] = '{32'hc2a14ef9};
test_output[3794] = '{32'h432cb739};
/*############ DEBUG ############
test_input[30352:30359] = '{89.3137327104, -29.0922515219, -17.6338773989, -60.2613973583, 11.2919179951, 91.9952531422, -16.6879311872, -80.6542428322};
test_label[3794] = '{-80.6542428322};
test_output[3794] = '{172.715713386};
############ END DEBUG ############*/
test_input[30360:30367] = '{32'h4277dafd, 32'hc1a320c2, 32'h428c617b, 32'hc02745fe, 32'hc245dd33, 32'h42ac77cd, 32'h421b7375, 32'hc2c22149};
test_label[3795] = '{32'h42ac77cd};
test_output[3795] = '{32'h33e76bfc};
/*############ DEBUG ############
test_input[30360:30367] = '{61.9638561514, -20.3909951271, 70.1903945393, -2.6136469376, -49.4660144138, 86.2339824188, 38.8627504538, -97.0650087351};
test_label[3795] = '{86.2339824188};
test_output[3795] = '{1.07764180835e-07};
############ END DEBUG ############*/
test_input[30368:30375] = '{32'hc2c7704c, 32'hc2958873, 32'h42c1f921, 32'h40a6771f, 32'h41ec592d, 32'hc166597c, 32'h418e6230, 32'hc18cca83};
test_label[3796] = '{32'hc2c7704c};
test_output[3796] = '{32'h4344b4b6};
/*############ DEBUG ############
test_input[30368:30375] = '{-99.7193284984, -74.7665034719, 96.9865787714, 5.20204092317, 29.5435427666, -14.3968467573, 17.7979422677, -17.5988817539};
test_label[3796] = '{-99.7193284984};
test_output[3796] = '{196.70590727};
############ END DEBUG ############*/
test_input[30376:30383] = '{32'h3ee01513, 32'h423925f2, 32'h41603478, 32'hc2c4f228, 32'hc2824223, 32'hc283b7aa, 32'hc203db09, 32'hc19d6a39};
test_label[3797] = '{32'hc19d6a39};
test_output[3797] = '{32'h4283ed87};
/*############ DEBUG ############
test_input[30376:30383] = '{0.437660781422, 46.2870558318, 14.0128101672, -98.4729590353, -65.1291696858, -65.8587187129, -32.9639023396, -19.6768674622};
test_label[3797] = '{-19.6768674622};
test_output[3797] = '{65.963923294};
############ END DEBUG ############*/
test_input[30384:30391] = '{32'h4014cc16, 32'hc2c45ce1, 32'hc243c347, 32'h41a2432d, 32'h42677f11, 32'hc21d8ab7, 32'hc103688d, 32'h41452980};
test_label[3798] = '{32'hc103688d};
test_output[3798] = '{32'h42842c9a};
/*############ DEBUG ############
test_input[30384:30391] = '{2.32495642596, -98.1814033327, -48.9407008145, 20.2828014028, 57.8740877473, -39.3854644866, -8.21302546166, 12.3226317609};
test_label[3798] = '{-8.21302546166};
test_output[3798] = '{66.087113209};
############ END DEBUG ############*/
test_input[30392:30399] = '{32'h429b7180, 32'hc24fa165, 32'hc242bfc6, 32'hc203e51a, 32'hc2582203, 32'hc271601d, 32'hc2c15272, 32'hc114d2c5};
test_label[3799] = '{32'hc242bfc6};
test_output[3799] = '{32'h42fcd164};
/*############ DEBUG ############
test_input[30392:30399] = '{77.7216832457, -51.9076104664, -48.6872790194, -32.9737302716, -54.0332159953, -60.3438602758, -96.6610281716, -9.30145705251};
test_label[3799] = '{-48.6872790194};
test_output[3799] = '{126.408962265};
############ END DEBUG ############*/
test_input[30400:30407] = '{32'hc1b81e4d, 32'h429fc38a, 32'h42aef5aa, 32'hc1f6cd56, 32'hc2bfb03b, 32'h427b1867, 32'h412022d6, 32'h4215b0c9};
test_label[3800] = '{32'hc2bfb03b};
test_output[3800] = '{32'h43375313};
/*############ DEBUG ############
test_input[30400:30407] = '{-23.0147958004, 79.881914288, 87.4798090033, -30.8502608022, -95.8441994009, 62.7738305504, 10.0085047684, 37.4226418349};
test_label[3800] = '{-95.8441994009};
test_output[3800] = '{183.324509785};
############ END DEBUG ############*/
test_input[30408:30415] = '{32'h42993669, 32'hc2ac4588, 32'h42902c2f, 32'hc10dd325, 32'hc25f8b61, 32'hc2b8dc7d, 32'h426c58d7, 32'h40b41cde};
test_label[3801] = '{32'h426c58d7};
test_output[3801] = '{32'h418c3e25};
/*############ DEBUG ############
test_input[30408:30415] = '{76.6062718714, -86.1358031966, 72.0862992094, -8.86404905835, -55.8861105547, -92.4306443656, 59.0867585502, 5.62852405533};
test_label[3801] = '{59.0867585502};
test_output[3801] = '{17.5303438052};
############ END DEBUG ############*/
test_input[30416:30423] = '{32'hc275affd, 32'hc220a4ec, 32'hc2b6c751, 32'hc21e4db9, 32'h42b818b7, 32'h41be9128, 32'hc2c6e770, 32'hc104b3bb};
test_label[3802] = '{32'hc2b6c751};
test_output[3802] = '{32'h43377004};
/*############ DEBUG ############
test_input[30416:30423] = '{-61.4218627007, -40.1610565401, -91.3892904624, -39.5759021933, 92.0482684141, 23.8208762894, -99.4520255205, -8.29387911869};
test_label[3802] = '{-91.3892904624};
test_output[3802] = '{183.437558877};
############ END DEBUG ############*/
test_input[30424:30431] = '{32'h420e3040, 32'hc2479049, 32'h416ced8d, 32'hc299b763, 32'h42499379, 32'hc1205d0c, 32'h42915f1c, 32'h420ab374};
test_label[3803] = '{32'hc1205d0c};
test_output[3803] = '{32'h42a56abd};
/*############ DEBUG ############
test_input[30424:30431] = '{35.547120286, -49.8909024778, 14.8079959327, -76.8581775308, 50.394017446, -10.0227161979, 72.6857600455, 34.6752457517};
test_label[3803] = '{-10.0227161979};
test_output[3803] = '{82.7084762436};
############ END DEBUG ############*/
test_input[30432:30439] = '{32'hc28734e5, 32'hc2c659cb, 32'h42608015, 32'h428e04cf, 32'hc19b21a5, 32'h42b3eddc, 32'hc2214785, 32'hc11eb63f};
test_label[3804] = '{32'h428e04cf};
test_output[3804] = '{32'h4197a434};
/*############ DEBUG ############
test_input[30432:30439] = '{-67.6033075202, -99.1753756347, 56.1250819816, 71.0093936823, -19.3914279942, 89.964570637, -40.3198428846, -9.91949341908};
test_label[3804] = '{71.0093936823};
test_output[3804] = '{18.9551769606};
############ END DEBUG ############*/
test_input[30440:30447] = '{32'hc146bf7e, 32'h42c3ccf6, 32'h429e3888, 32'h429b674e, 32'hc1cf9b9d, 32'hc26d3745, 32'h424fe3dd, 32'h42927b10};
test_label[3805] = '{32'h429b674e};
test_output[3805] = '{32'h41a196a1};
/*############ DEBUG ############
test_input[30440:30447] = '{-12.4217512449, 97.900313434, 79.1104162596, 77.7017640041, -25.9509825179, -59.3039752972, 51.9725226398, 73.2403569978};
test_label[3805] = '{77.7017640041};
test_output[3805] = '{20.1985494385};
############ END DEBUG ############*/
test_input[30448:30455] = '{32'h42243f0a, 32'h42084649, 32'hc1c05579, 32'hc2adab42, 32'hc27da744, 32'h428e1384, 32'h42080de1, 32'hc13faa4e};
test_label[3806] = '{32'h42243f0a};
test_output[3806] = '{32'h41efcffb};
/*############ DEBUG ############
test_input[30448:30455] = '{41.0615602022, 34.0686383431, -24.0417345277, -86.8344870005, -63.4133452386, 71.0381137364, 34.0135517498, -11.9790779474};
test_label[3806] = '{41.0615602022};
test_output[3806] = '{29.9765535343};
############ END DEBUG ############*/
test_input[30456:30463] = '{32'hc22f618d, 32'hc2852656, 32'hc0c1debc, 32'h4258ecb4, 32'hc1ade8ff, 32'hc28b7348, 32'h3f168466, 32'hc245f7e9};
test_label[3807] = '{32'hc0c1debc};
test_output[3807] = '{32'h4271288b};
/*############ DEBUG ############
test_input[30456:30463] = '{-43.8452640249, -66.5748758926, -6.05843945927, 54.2311545565, -21.7387668664, -69.7251580902, 0.587957749627, -49.4921005181};
test_label[3807] = '{-6.05843945927};
test_output[3807] = '{60.2895940158};
############ END DEBUG ############*/
test_input[30464:30471] = '{32'h42b716dc, 32'hc223901f, 32'hc2a82d56, 32'hc2b85e70, 32'h429d164b, 32'hc2c6f7a5, 32'hc2b05c66, 32'h42a04494};
test_label[3808] = '{32'hc223901f};
test_output[3808] = '{32'h43046f76};
/*############ DEBUG ############
test_input[30464:30471] = '{91.5446450627, -40.8907431862, -84.0885503822, -92.184445069, 78.5435432966, -99.4836825113, -88.18046324, 80.1339429019};
test_label[3808] = '{-40.8907431862};
test_output[3808] = '{132.435401583};
############ END DEBUG ############*/
test_input[30472:30479] = '{32'h42b33038, 32'h42a1e3c0, 32'h41da4557, 32'h42b5d59f, 32'hc2a30d9d, 32'h42affa92, 32'hc1b3a07c, 32'hc1b37dbf};
test_label[3809] = '{32'h42b33038};
test_output[3809] = '{32'h3fcce044};
/*############ DEBUG ############
test_input[30472:30479] = '{89.5941777967, 80.9448225817, 27.2838581341, 90.9172306971, -81.526585476, 87.9893947189, -22.4533615068, -22.4363989751};
test_label[3809] = '{89.5941777967};
test_output[3809] = '{1.6005940221};
############ END DEBUG ############*/
test_input[30480:30487] = '{32'h42af8341, 32'h422511ea, 32'h42657629, 32'h4258f0b7, 32'h41e6bbbd, 32'hc2808d13, 32'h41f1a83d, 32'hc10d83fd};
test_label[3810] = '{32'h41e6bbbd};
test_output[3810] = '{32'h426ba8a3};
/*############ DEBUG ############
test_input[30480:30487] = '{87.7563542802, 41.2674935939, 57.3653925053, 54.2350722808, 28.8416684817, -64.2755375374, 30.2071476633, -8.84472347147};
test_label[3810] = '{28.8416684817};
test_output[3810] = '{58.9146857985};
############ END DEBUG ############*/
test_input[30488:30495] = '{32'h42aea311, 32'h4264249d, 32'h425d4a2c, 32'h42c5de2f, 32'h421f259f, 32'hc2c65fa9, 32'h42bf36ac, 32'h42826427};
test_label[3811] = '{32'h42bf36ac};
test_output[3811] = '{32'h40573235};
/*############ DEBUG ############
test_input[30488:30495] = '{87.3184864005, 57.0357539898, 55.3224333384, 98.933949755, 39.786740427, -99.1868325763, 95.6067846255, 65.1956112711};
test_label[3811] = '{95.6067846255};
test_output[3811] = '{3.36243935713};
############ END DEBUG ############*/
test_input[30496:30503] = '{32'hc24e9dfa, 32'h4253e6ae, 32'h4233d25b, 32'hc18d4599, 32'hc25a3aa6, 32'h429eaf29, 32'h42a323ec, 32'hc2057bba};
test_label[3812] = '{32'hc2057bba};
test_output[3812] = '{32'h42e6162d};
/*############ DEBUG ############
test_input[30496:30503] = '{-51.6542757179, 52.9752749696, 44.9554238262, -17.6589837151, -54.5572730308, 79.342107291, 81.5701619286, -33.3708282303};
test_label[3812] = '{-33.3708282303};
test_output[3812] = '{115.043310091};
############ END DEBUG ############*/
test_input[30504:30511] = '{32'hc2840015, 32'h41f37337, 32'h41034d56, 32'hc28ff357, 32'hc24deec7, 32'hc23a3c33, 32'h41563ec0, 32'h429e129c};
test_label[3813] = '{32'h41f37337};
test_output[3813] = '{32'h42426b9d};
/*############ DEBUG ############
test_input[30504:30511] = '{-66.0001623814, 30.4312564542, 8.20638079649, -71.9752699043, -51.4831812359, -46.5587891806, 13.3903202078, 79.0363467657};
test_label[3813] = '{30.4312564542};
test_output[3813] = '{48.6050903115};
############ END DEBUG ############*/
test_input[30512:30519] = '{32'hc1a748ed, 32'h3f65db99, 32'hc2a1b189, 32'h4233aefd, 32'hc2742acd, 32'h42c5c667, 32'h424e9aec, 32'h42b2efca};
test_label[3814] = '{32'h4233aefd};
test_output[3814] = '{32'h4257dde6};
/*############ DEBUG ############
test_input[30512:30519] = '{-20.9106079458, 0.897882039839, -80.8467463023, 44.9208871572, -61.0417957992, 98.8875023742, 51.6512900547, 89.4683366097};
test_label[3814] = '{44.9208871572};
test_output[3814] = '{53.9666963674};
############ END DEBUG ############*/
test_input[30520:30527] = '{32'h4226119a, 32'hc2b2204e, 32'hc2b92e37, 32'hc28d36e8, 32'h41800879, 32'h418296ec, 32'hc1eb7bba, 32'h40d1a225};
test_label[3815] = '{32'h41800879};
test_output[3815] = '{32'h41cc1abc};
/*############ DEBUG ############
test_input[30520:30527] = '{41.5171908096, -89.0630954589, -92.5902654494, -70.6072374845, 16.0041362361, 16.3236918321, -29.4354128931, 6.55104293589};
test_label[3815] = '{16.0041362361};
test_output[3815] = '{25.5130545735};
############ END DEBUG ############*/
test_input[30528:30535] = '{32'h42983549, 32'hc2743104, 32'h42c197ef, 32'h42c46515, 32'hc20a6cc5, 32'h42c40c1b, 32'hc2836226, 32'hc2788f8b};
test_label[3816] = '{32'h42983549};
test_output[3816] = '{32'h41b6a1df};
/*############ DEBUG ############
test_input[30528:30535] = '{76.104073701, -61.0478665229, 96.7967432372, 98.1974285068, -34.6062189897, 98.0236467004, -65.6916931284, -62.1401776537};
test_label[3816] = '{76.104073701};
test_output[3816] = '{22.8290384951};
############ END DEBUG ############*/
test_input[30536:30543] = '{32'hc29006ed, 32'hc1d3606b, 32'h41bbbaea, 32'h42194d64, 32'h41f6e670, 32'hc2a7381f, 32'hc2947ff9, 32'hc2871d23};
test_label[3817] = '{32'hc2a7381f};
test_output[3817] = '{32'h42f3df1c};
/*############ DEBUG ############
test_input[30536:30543] = '{-72.0135246429, -26.4220799586, 23.4662660379, 38.3255765272, 30.8625186415, -83.6096109976, -74.2499431025, -67.5569055955};
test_label[3817] = '{-83.6096109976};
test_output[3817] = '{121.935761611};
############ END DEBUG ############*/
test_input[30544:30551] = '{32'hc2a38210, 32'hc243076d, 32'h42548af8, 32'h410056ee, 32'hc1f3367f, 32'h426d2750, 32'h40abf017, 32'h42b92287};
test_label[3818] = '{32'h42b92287};
test_output[3818] = '{32'h27780000};
/*############ DEBUG ############
test_input[30544:30551] = '{-81.7540305473, -48.7572513862, 53.1357126564, 8.02122327255, -30.4016088877, 59.2883906318, 5.37305789408, 92.5674356247};
test_label[3818] = '{92.5674356247};
test_output[3818] = '{3.44169137634e-15};
############ END DEBUG ############*/
test_input[30552:30559] = '{32'h42a45acb, 32'hc19134ee, 32'h41a3d58b, 32'hc1fa609b, 32'hc29ac767, 32'h40dfa913, 32'hc18ca997, 32'h42acd1e8};
test_label[3819] = '{32'hc29ac767};
test_output[3819] = '{32'h4323d058};
/*############ DEBUG ############
test_input[30552:30559] = '{82.177328769, -18.1508450598, 20.4792697814, -31.29717154, -77.3894555446, 6.98938876966, -17.5828066295, 86.4099759583};
test_label[3819] = '{-77.3894555446};
test_output[3819] = '{163.813841103};
############ END DEBUG ############*/
test_input[30560:30567] = '{32'hc1b0df01, 32'h409d7163, 32'h42b2f233, 32'hc2878c3d, 32'hc0fe9ee3, 32'h4221972b, 32'h42286ea7, 32'hc2c25ff7};
test_label[3820] = '{32'hc2878c3d};
test_output[3820] = '{32'h431d3f38};
/*############ DEBUG ############
test_input[30560:30567] = '{-22.1088883714, 4.92009109192, 89.4730437012, -67.7738995495, -7.95689527985, 40.3976261066, 42.108057963, -97.1874327171};
test_label[3820] = '{-67.7738995495};
test_output[3820] = '{157.246943251};
############ END DEBUG ############*/
test_input[30568:30575] = '{32'hc2c1a354, 32'h40d681f5, 32'hc0a5b911, 32'hc27a45fa, 32'h4299b033, 32'h405cc580, 32'hc283742c, 32'hc2af7133};
test_label[3821] = '{32'hc0a5b911};
test_output[3821] = '{32'h42a40bc4};
/*############ DEBUG ############
test_input[30568:30575] = '{-96.8189978107, 6.70336367613, -5.17884103519, -62.5683363978, 76.8441367164, 3.44955455601, -65.7268958587, -87.7210947321};
test_label[3821] = '{-5.17884103519};
test_output[3821] = '{82.0229777516};
############ END DEBUG ############*/
test_input[30576:30583] = '{32'hc25cc842, 32'h42b85929, 32'h413fef1c, 32'h42378c06, 32'hc10afe25, 32'h428a53eb, 32'h410daf51, 32'hc1ae0c05};
test_label[3822] = '{32'h42378c06};
test_output[3822] = '{32'h4239264b};
/*############ DEBUG ############
test_input[30576:30583] = '{-55.1955648887, 92.1741385039, 11.9958760481, 45.8867415746, -8.68704695808, 69.1639036141, 8.85530173435, -21.7558690774};
test_label[3822] = '{45.8867415746};
test_output[3822] = '{46.2873969294};
############ END DEBUG ############*/
test_input[30584:30591] = '{32'h428e5030, 32'hc15ef776, 32'hc28b0edb, 32'h3fcc8125, 32'h42c28e45, 32'h4281a0d4, 32'h428ae268, 32'hc296facd};
test_label[3823] = '{32'h428ae268};
test_output[3823] = '{32'h41deaf75};
/*############ DEBUG ############
test_input[30584:30591] = '{71.1566143905, -13.935415223, -69.5290129523, 1.59769117772, 97.2778705028, 64.8141183859, 69.4421975133, -75.4898455438};
test_label[3823] = '{69.4421975133};
test_output[3823] = '{27.8356729896};
############ END DEBUG ############*/
test_input[30592:30599] = '{32'h42646083, 32'h4215112b, 32'hc2bb00ac, 32'h4293347c, 32'hc265541a, 32'hc250052a, 32'hc2b5b220, 32'h42c59c1a};
test_label[3824] = '{32'h4293347c};
test_output[3824] = '{32'h41c99e76};
/*############ DEBUG ############
test_input[30592:30599] = '{57.0942489096, 37.2667661254, -93.5013084717, 73.602509048, -57.3321300694, -52.0050429296, -90.8479033556, 98.804882366};
test_label[3824] = '{73.602509048};
test_output[3824] = '{25.202373318};
############ END DEBUG ############*/
test_input[30600:30607] = '{32'hc2b41834, 32'hc205ec7a, 32'hc1165b5d, 32'hc29b92c9, 32'h42832416, 32'hc2b44f84, 32'hc21b36e2, 32'hc16abf2c};
test_label[3825] = '{32'hc21b36e2};
test_output[3825] = '{32'h42d0bf88};
/*############ DEBUG ############
test_input[30600:30607] = '{-90.0472692912, -33.4809328977, -9.39730545944, -77.7866931057, 65.5704831946, -90.1553070846, -38.8035981084, -14.6716726118};
test_label[3825] = '{-38.8035981084};
test_output[3825] = '{104.374081303};
############ END DEBUG ############*/
test_input[30608:30615] = '{32'h428998a5, 32'h3f72caa0, 32'h422c6f8b, 32'h42b0619a, 32'h40c4ab07, 32'hc2baa1ba, 32'hc173487d, 32'hc230dfff};
test_label[3826] = '{32'hc2baa1ba};
test_output[3826] = '{32'h433581aa};
/*############ DEBUG ############
test_input[30608:30615] = '{68.798136691, 0.948404285564, 43.1089294149, 88.1906289385, 6.14587754497, -93.3158693424, -15.205196924, -44.2187443718};
test_label[3826] = '{-93.3158693424};
test_output[3826] = '{181.506498285};
############ END DEBUG ############*/
test_input[30616:30623] = '{32'h4276af56, 32'h42a4576d, 32'hc2900a04, 32'hc1cec73c, 32'h42220de3, 32'hc2aecf1a, 32'hc2b0fb06, 32'h428c0e56};
test_label[3827] = '{32'hc2900a04};
test_output[3827] = '{32'h431a30b9};
/*############ DEBUG ############
test_input[30616:30623] = '{61.6712279345, 82.1707516261, -72.0195594117, -25.8472827, 40.5135626281, -87.4044915695, -88.4902831072, 70.0279988663};
test_label[3827] = '{-72.0195594117};
test_output[3827] = '{154.190316366};
############ END DEBUG ############*/
test_input[30624:30631] = '{32'hc075d706, 32'h42bf1aca, 32'h42c7f83c, 32'h426090b2, 32'h416f828c, 32'h41feb389, 32'hc0fb72f2, 32'hc29771cc};
test_label[3828] = '{32'hc0fb72f2};
test_output[3828] = '{32'h42d7b577};
/*############ DEBUG ############
test_input[30624:30631] = '{-3.84124890646, 95.552326, 99.9848292263, 56.1413040887, 14.9693719925, 31.8376634805, -7.85778127459, -75.7222614328};
test_label[3828] = '{-7.85778127459};
test_output[3828] = '{107.854425135};
############ END DEBUG ############*/
test_input[30632:30639] = '{32'h3e22bb30, 32'h423c5dce, 32'hc25c1126, 32'hc2288d24, 32'h42bc45ec, 32'h412c271c, 32'hc267dc76, 32'h42993837};
test_label[3829] = '{32'hc25c1126};
test_output[3829] = '{32'h4315273f};
/*############ DEBUG ############
test_input[30632:30639] = '{0.158917195237, 47.0916077014, -55.0167454373, -42.1378315514, 94.1365665605, 10.7595486126, -57.9652934748, 76.6097957555};
test_label[3829] = '{-55.0167454373};
test_output[3829] = '{149.153312022};
############ END DEBUG ############*/
test_input[30640:30647] = '{32'h426056bc, 32'h429df3af, 32'hc20120a1, 32'hc1aa6270, 32'hc2a6e9f9, 32'h42b3de45, 32'h425ab88e, 32'h412bd210};
test_label[3830] = '{32'hc1aa6270};
test_output[3830] = '{32'h42de76e3};
/*############ DEBUG ############
test_input[30640:30647] = '{56.0847028734, 78.9759418432, -32.2818657476, -21.2980657027, -83.4569757401, 89.9341177695, 54.6802286579, 10.7387847266};
test_label[3830] = '{-21.2980657027};
test_output[3830] = '{111.232200887};
############ END DEBUG ############*/
test_input[30648:30655] = '{32'hc219d70d, 32'hc19b48fd, 32'h42b6ed82, 32'hc1ea92d8, 32'hc2998238, 32'hc2aca182, 32'h4247c988, 32'hc19e78d1};
test_label[3831] = '{32'h42b6ed82};
test_output[3831] = '{32'h80000000};
/*############ DEBUG ############
test_input[30648:30655] = '{-38.4600103687, -19.4106394006, 91.4638848754, -29.3217008594, -76.7543366385, -86.3154461101, 49.9468068014, -19.8089925391};
test_label[3831] = '{91.4638848754};
test_output[3831] = '{-0.0};
############ END DEBUG ############*/
test_input[30656:30663] = '{32'h4298fb4e, 32'hc29ab966, 32'hc25d2449, 32'h40ff294d, 32'h42b10638, 32'hc2135012, 32'h4255cde4, 32'hc290144f};
test_label[3832] = '{32'h40ff294d};
test_output[3832] = '{32'h42a113a4};
/*############ DEBUG ############
test_input[30656:30663] = '{76.4908312726, -77.362106953, -55.2854358786, 7.97379179348, 88.5121493871, -36.8281952363, 53.4510667315, -72.0396687659};
test_label[3832] = '{7.97379179348};
test_output[3832] = '{80.5383636082};
############ END DEBUG ############*/
test_input[30664:30671] = '{32'h4236e6b3, 32'hbf61b84c, 32'h41f16bb7, 32'hc21b761b, 32'h42bf9800, 32'h4228d4be, 32'h42458f36, 32'hbf410d16};
test_label[3833] = '{32'hbf61b84c};
test_output[3833] = '{32'h42c15b71};
/*############ DEBUG ############
test_input[30664:30671] = '{45.7252910563, -0.881718417825, 30.1775951333, -38.8653373389, 95.7968781102, 42.2077554219, 49.3898533644, -0.754105941547};
test_label[3833] = '{-0.881718417825};
test_output[3833] = '{96.678596528};
############ END DEBUG ############*/
test_input[30672:30679] = '{32'hc1af0594, 32'hc29d6f4b, 32'h42a35561, 32'hc1e8d235, 32'h429d06b5, 32'hc049c8ca, 32'h428fec79, 32'hc23544be};
test_label[3834] = '{32'h42a35561};
test_output[3834] = '{32'h3d2b7d7c};
/*############ DEBUG ############
test_input[30672:30679] = '{-21.8777233107, -78.7173727815, 81.6667584998, -29.102639703, 78.513097908, -3.15288030937, 71.9618637473, -45.3171309064};
test_label[3834] = '{81.6667584998};
test_output[3834] = '{0.0418677199483};
############ END DEBUG ############*/
test_input[30680:30687] = '{32'h3f41bb5e, 32'h42906f75, 32'h42a79878, 32'hc2bc2d95, 32'h41bf2e09, 32'hc2a72d87, 32'hc1ea3187, 32'hc10655e8};
test_label[3835] = '{32'hc2bc2d95};
test_output[3835] = '{32'h4331e307};
/*############ DEBUG ############
test_input[30680:30687] = '{0.756765252153, 72.2176881907, 83.7977896412, -94.0890270282, 23.8974778094, -83.5889230414, -29.274183387, -8.39597286548};
test_label[3835] = '{-94.0890270282};
test_output[3835] = '{177.88682602};
############ END DEBUG ############*/
test_input[30688:30695] = '{32'hc010c6bf, 32'hc2b83c24, 32'hc275fa4c, 32'hc2beab64, 32'hc18b7e33, 32'hc23bebdf, 32'hc1fd5b10, 32'h41919afc};
test_label[3836] = '{32'hc2beab64};
test_output[3836] = '{32'h42e31223};
/*############ DEBUG ############
test_input[30688:30695] = '{-2.26213048835, -92.1174642495, -61.4944305105, -95.3347506157, -17.4366197705, -46.980342676, -31.6694649902, 18.2006756722};
test_label[3836] = '{-95.3347506157};
test_output[3836] = '{113.535426289};
############ END DEBUG ############*/
test_input[30696:30703] = '{32'h427dd975, 32'h422548ca, 32'hc283b01e, 32'hc2b85223, 32'h423cb083, 32'h42b21e78, 32'h414ea6ef, 32'h42b563c1};
test_label[3837] = '{32'hc2b85223};
test_output[3837] = '{32'h43370887};
/*############ DEBUG ############
test_input[30696:30703] = '{63.4623622795, 41.3210849584, -65.8439756397, -92.1604248439, 47.1723758941, 89.0595056639, 12.9157549646, 90.6948350953};
test_label[3837] = '{-92.1604248439};
test_output[3837] = '{183.033312529};
############ END DEBUG ############*/
test_input[30704:30711] = '{32'h42c4d5e8, 32'hc2316284, 32'hc22585c0, 32'hc2a63a1d, 32'hc1618169, 32'hc029bf8b, 32'hc2878230, 32'hc1f97533};
test_label[3838] = '{32'hc029bf8b};
test_output[3838] = '{32'h42ca23e4};
/*############ DEBUG ############
test_input[30704:30711] = '{98.4177861158, -44.3462083183, -41.3806151245, -83.1135007143, -14.094094263, -2.65231585842, -67.7542692448, -31.1822264276};
test_label[3838] = '{-2.65231585842};
test_output[3838] = '{101.070101974};
############ END DEBUG ############*/
test_input[30712:30719] = '{32'hc22ee508, 32'h42c7f68d, 32'hc2195317, 32'h422882c9, 32'h410c825c, 32'h4247154e, 32'hc20fc908, 32'h428d0621};
test_label[3839] = '{32'h42c7f68d};
test_output[3839] = '{32'h2a332000};
/*############ DEBUG ############
test_input[30712:30719] = '{-43.7236638195, 99.9815454141, -38.3311437189, 42.1277215352, 8.78182606865, 49.7708066462, -35.9463204926, 70.5119667853};
test_label[3839] = '{99.9815454141};
test_output[3839] = '{1.59094959429e-13};
############ END DEBUG ############*/
test_input[30720:30727] = '{32'h42971c0d, 32'h42a90e10, 32'hc245290a, 32'h41ef3f4a, 32'hc28979af, 32'h4246b7b6, 32'hc2a74460, 32'h4288a7d9};
test_label[3840] = '{32'h41ef3f4a};
test_output[3840] = '{32'h425a7c9c};
/*############ DEBUG ############
test_input[30720:30727] = '{75.5547883019, 84.5274643601, -49.2900777506, 29.9059026647, -68.7376641952, 49.679404707, -83.6335422302, 68.3278288435};
test_label[3840] = '{29.9059026647};
test_output[3840] = '{54.6216886078};
############ END DEBUG ############*/
test_input[30728:30735] = '{32'hc1da5da5, 32'h42c41762, 32'hc274bda7, 32'h425596d0, 32'hc1bb6378, 32'h416c2e3c, 32'hc2778e77, 32'h4229dbcd};
test_label[3841] = '{32'hc1bb6378};
test_output[3841] = '{32'h42f2f040};
/*############ DEBUG ############
test_input[30728:30735] = '{-27.2957247345, 98.0456686012, -61.1852080817, 53.3972777917, -23.4235684465, 14.7612879298, -61.8891239847, 42.4646475239};
test_label[3841] = '{-23.4235684465};
test_output[3841] = '{121.469237048};
############ END DEBUG ############*/
test_input[30736:30743] = '{32'h41bcf577, 32'hc213fe3a, 32'hc1f3a96c, 32'hc219b49d, 32'hc29fb7cc, 32'hc21d7c6b, 32'h42383ee5, 32'h41da1c30};
test_label[3842] = '{32'hc219b49d};
test_output[3842] = '{32'h42a8f9c1};
/*############ DEBUG ############
test_input[30736:30743] = '{23.6198565231, -36.998268319, -30.4577263674, -38.4263813317, -79.8589802424, -39.3715035062, 46.061421163, 27.2637627388};
test_label[3842] = '{-38.4263813317};
test_output[3842] = '{84.4878025017};
############ END DEBUG ############*/
test_input[30744:30751] = '{32'hc19092d1, 32'hc2070549, 32'hc141ce96, 32'h411e6291, 32'hc1fbd7de, 32'hc26c7dad, 32'hc1486d99, 32'hc1c100f7};
test_label[3843] = '{32'hc26c7dad};
test_output[3843] = '{32'h428a0b29};
/*############ DEBUG ############
test_input[30744:30751] = '{-18.0716880757, -33.7551615555, -12.1129363757, 9.89906414218, -31.4804046956, -59.1227301852, -12.5267576641, -24.1254711765};
test_label[3843] = '{-59.1227301852};
test_output[3843] = '{69.0217943278};
############ END DEBUG ############*/
test_input[30752:30759] = '{32'h419fb088, 32'hc1fcd732, 32'hc2c46e24, 32'hc26be56d, 32'h42ad37ba, 32'hc2ae41e9, 32'h423198c8, 32'h42314c09};
test_label[3844] = '{32'h419fb088};
test_output[3844] = '{32'h42854b98};
/*############ DEBUG ############
test_input[30752:30759] = '{19.9611967402, -31.6050757859, -98.2151174232, -58.9740483445, 86.6088419492, -87.1287271237, 44.3992004258, 44.3242528661};
test_label[3844] = '{19.9611967402};
test_output[3844] = '{66.6476452091};
############ END DEBUG ############*/
test_input[30760:30767] = '{32'h42282a80, 32'hc21b7e8e, 32'h4215eee6, 32'h412571db, 32'hc227dd55, 32'h415074ac, 32'h40d9af63, 32'h414d1707};
test_label[3845] = '{32'h42282a80};
test_output[3845] = '{32'h3c2ad31a};
/*############ DEBUG ############
test_input[30760:30767] = '{42.0415052186, -38.8735873005, 37.4832997596, 10.3402969029, -41.9661453488, 13.0284840151, 6.80265955672, 12.8181215716};
test_label[3845] = '{42.0415052186};
test_output[3845] = '{0.0104263070573};
############ END DEBUG ############*/
test_input[30768:30775] = '{32'hc1e0cad6, 32'h42318d33, 32'h41e22056, 32'h42837ff3, 32'h421b7e23, 32'h3fbcff9b, 32'hc1d5e4ad, 32'h41fa01bc};
test_label[3846] = '{32'h42837ff3};
test_output[3846] = '{32'h3011b552};
/*############ DEBUG ############
test_input[30768:30775] = '{-28.0990405606, 44.3878912151, 28.2657897749, 65.7498985026, 38.8731785586, 1.47655040366, -26.7366583672, 31.2508471814};
test_label[3846] = '{65.7498985026};
test_output[3846] = '{5.30083643787e-10};
############ END DEBUG ############*/
test_input[30776:30783] = '{32'h42bd1ffe, 32'h416e33fd, 32'h425081b5, 32'hc2545701, 32'h427508fc, 32'hc1fb231b, 32'h41da5abe, 32'h4289db4d};
test_label[3847] = '{32'h42bd1ffe};
test_output[3847] = '{32'h2d01a480};
/*############ DEBUG ############
test_input[30776:30783] = '{94.5624867212, 14.8876919834, 52.1266658145, -53.0849666255, 61.2587754736, -31.3921410499, 27.2943084945, 68.9283230381};
test_label[3847] = '{94.5624867212};
test_output[3847] = '{7.36932737058e-12};
############ END DEBUG ############*/
test_input[30784:30791] = '{32'hc23aa8ef, 32'hc21aaa2b, 32'hc2bc477e, 32'h41cda30e, 32'h42a5fdb9, 32'hc1416d73, 32'hc208bb54, 32'h42bc242f};
test_label[3848] = '{32'h42a5fdb9};
test_output[3848] = '{32'h413133c0};
/*############ DEBUG ############
test_input[30784:30791] = '{-46.6649733405, -38.6661803505, -94.1396347269, 25.7046157261, 82.9955554535, -12.0892212101, -34.1829371805, 94.070674241};
test_label[3848] = '{82.9955554535};
test_output[3848] = '{11.0751342804};
############ END DEBUG ############*/
test_input[30792:30799] = '{32'h41b53891, 32'hc2841869, 32'hc2bb4eb4, 32'h4151d60b, 32'hc2992c3d, 32'hc09c8e22, 32'hc28d4b86, 32'h42b3c1a2};
test_label[3849] = '{32'h42b3c1a2};
test_output[3849] = '{32'h80000000};
/*############ DEBUG ############
test_input[30792:30799] = '{22.6526203144, -66.0476723035, -93.6537167556, 13.1147565544, -76.5864036202, -4.89235024651, -70.6475056067, 89.8781854091};
test_label[3849] = '{89.8781854091};
test_output[3849] = '{-0.0};
############ END DEBUG ############*/
test_input[30800:30807] = '{32'hc262a9ab, 32'h4271ae9d, 32'hc21d48ae, 32'h42c69ecb, 32'hc232ddc2, 32'hc289b881, 32'h41971e7b, 32'h4203aba1};
test_label[3850] = '{32'hc289b881};
test_output[3850] = '{32'h43282ba6};
/*############ DEBUG ############
test_input[30800:30807] = '{-56.6656908248, 60.4205221085, -39.3209758473, 99.3101430346, -44.7165593598, -68.8603616142, 18.8898836996, 32.9176049305};
test_label[3850] = '{-68.8603616142};
test_output[3850] = '{168.170504649};
############ END DEBUG ############*/
test_input[30808:30815] = '{32'h414af9e5, 32'hc28fa398, 32'h40f4644d, 32'hc239e013, 32'hc24dd011, 32'h4274c60f, 32'h42964968, 32'hc28c00c8};
test_label[3851] = '{32'hc28c00c8};
test_output[3851] = '{32'h43112518};
/*############ DEBUG ############
test_input[30808:30815] = '{12.6860095249, -71.8195172184, 7.63724387141, -46.468821156, -51.453189367, 61.1934179272, 75.1433734115, -70.0015278563};
test_label[3851] = '{-70.0015278563};
test_output[3851] = '{145.144902142};
############ END DEBUG ############*/
test_input[30816:30823] = '{32'h41bf263c, 32'h414f70cf, 32'hc210dae9, 32'hc224cb46, 32'h425844f8, 32'hc2aebf28, 32'h41485eea, 32'hc298c0a3};
test_label[3852] = '{32'h41bf263c};
test_output[3852] = '{32'h41f163b4};
/*############ DEBUG ############
test_input[30816:30823] = '{23.8936691378, 12.9650415519, -36.2137780484, -41.198510987, 54.0673513854, -87.3733544531, 12.5231723463, -76.376244498};
test_label[3852] = '{23.8936691378};
test_output[3852] = '{30.1736822476};
############ END DEBUG ############*/
test_input[30824:30831] = '{32'hc2149f5e, 32'h42ae07b1, 32'h41d869e9, 32'h429e74ae, 32'hc23ef156, 32'hc24f43c5, 32'hc1d35757, 32'hc14cbd11};
test_label[3853] = '{32'h429e74ae};
test_output[3853] = '{32'h40f9339b};
/*############ DEBUG ############
test_input[30824:30831] = '{-37.1556332777, 87.0150225576, 27.0517131149, 79.227887884, -47.7356806484, -51.8161830561, -26.41764731, -12.7961588732};
test_label[3853] = '{79.227887884};
test_output[3853] = '{7.78754962791};
############ END DEBUG ############*/
test_input[30832:30839] = '{32'hc22052db, 32'hc2160faa, 32'hc2398c53, 32'hc1cb0116, 32'hc25748c7, 32'hc20ffa83, 32'h42b39f0e, 32'hc29abc41};
test_label[3854] = '{32'hc22052db};
test_output[3854] = '{32'h4301e43e};
/*############ DEBUG ############
test_input[30832:30839] = '{-40.0809129834, -37.5152978715, -46.3870358558, -25.3755309154, -53.8210732725, -35.9946415214, 89.8106556749, -77.3676858696};
test_label[3854] = '{-40.0809129834};
test_output[3854] = '{129.891568658};
############ END DEBUG ############*/
test_input[30840:30847] = '{32'hc2a63c4f, 32'hc191323e, 32'hc25042ae, 32'hc2909012, 32'hc26e49e5, 32'hc264feb1, 32'hc1fe96e8, 32'hc2374c03};
test_label[3855] = '{32'hc1fe96e8};
test_output[3855] = '{32'h415ac957};
/*############ DEBUG ############
test_input[30840:30847] = '{-83.1177931251, -18.1495314283, -52.0651156896, -72.2813892113, -59.5721612247, -57.2487209565, -31.8236851246, -45.8242302624};
test_label[3855] = '{-31.8236851246};
test_output[3855] = '{13.6741548482};
############ END DEBUG ############*/
test_input[30848:30855] = '{32'hc1f3b77a, 32'hc242f1c6, 32'h41262e5e, 32'h4224d1c3, 32'hc228a6d8, 32'h41896f73, 32'hc22b4ddf, 32'hc215b916};
test_label[3856] = '{32'hc22b4ddf};
test_output[3856] = '{32'h42a80fd1};
/*############ DEBUG ############
test_input[30848:30855] = '{-30.4645889625, -48.7361061887, 10.3863204794, 41.2048451828, -42.1629344393, 17.1794191332, -42.8260452651, -37.4307471865};
test_label[3856] = '{-42.8260452651};
test_output[3856] = '{84.030890448};
############ END DEBUG ############*/
test_input[30856:30863] = '{32'hc25e8254, 32'h4285fe76, 32'hbcd0814a, 32'hc183f069, 32'h42a63017, 32'h423b6a5e, 32'hc22c4ad9, 32'h4134faee};
test_label[3857] = '{32'hc25e8254};
test_output[3857] = '{32'h430ab8a1};
/*############ DEBUG ############
test_input[30856:30863] = '{-55.6272753841, 66.9969926921, -0.0254522746562, -16.4923873893, 83.0939244687, 46.8538740588, -43.0730934666, 11.3112619184};
test_label[3857] = '{-55.6272753841};
test_output[3857] = '{138.721199955};
############ END DEBUG ############*/
test_input[30864:30871] = '{32'hc2638913, 32'h42c1fbc9, 32'h4263c392, 32'hc19e3729, 32'hc14896eb, 32'hc283bb8b, 32'h41e9ce50, 32'h41f547ba};
test_label[3858] = '{32'h41e9ce50};
test_output[3858] = '{32'h42878835};
/*############ DEBUG ############
test_input[30864:30871] = '{-56.8838610115, 96.9917665889, 56.9409885379, -19.7769339634, -12.5368447978, -65.8662924571, 29.2257377799, 30.6600235357};
test_label[3858] = '{29.2257377799};
test_output[3858] = '{67.766028809};
############ END DEBUG ############*/
test_input[30872:30879] = '{32'hc22a9fd1, 32'hc283b4e3, 32'hc22c5cc1, 32'h4238b04c, 32'h40af59e2, 32'h42b2670e, 32'h42a9fd3e, 32'h427ecb6e};
test_label[3859] = '{32'h427ecb6e};
test_output[3859] = '{32'h41cc23a3};
/*############ DEBUG ############
test_input[30872:30879] = '{-42.6560698821, -65.8532909025, -43.0905800336, 46.1721665573, 5.47972185409, 89.2012756637, 84.9946132654, 63.6986604219};
test_label[3859] = '{63.6986604219};
test_output[3859] = '{25.5174013884};
############ END DEBUG ############*/
test_input[30880:30887] = '{32'h4178158e, 32'hc2306eca, 32'hc2b3dc1f, 32'h4283fe5c, 32'h42b72cfb, 32'h42aa802f, 32'h41bffd7b, 32'h4263fb0d};
test_label[3860] = '{32'hc2b3dc1f};
test_output[3860] = '{32'h43358501};
/*############ DEBUG ############
test_input[30880:30887] = '{15.5052623375, -44.1081937521, -89.9299207719, 65.9967991096, 91.5878544292, 85.2503598122, 23.9987698104, 56.9951655361};
test_label[3860] = '{-89.9299207719};
test_output[3860] = '{181.519542367};
############ END DEBUG ############*/
test_input[30888:30895] = '{32'hc2a2dada, 32'hc1b881f8, 32'h426e9cb4, 32'hc0d755b6, 32'hc216bc94, 32'hc23ae596, 32'h42b8f041, 32'h426c9960};
test_label[3861] = '{32'hc23ae596};
test_output[3861] = '{32'h430b3186};
/*############ DEBUG ############
test_input[30888:30895] = '{-81.4274460592, -23.0634605759, 59.6530316173, -6.72921289846, -37.6841573032, -46.7242068855, 92.4692459024, 59.1497819197};
test_label[3861] = '{-46.7242068855};
test_output[3861] = '{139.193452788};
############ END DEBUG ############*/
test_input[30896:30903] = '{32'hc26cd170, 32'h4284e8ae, 32'h408c3498, 32'hc24637f2, 32'hc267d8a0, 32'h42aa74a2, 32'h428434a4, 32'hc1c306b8};
test_label[3862] = '{32'h42aa74a2};
test_output[3862] = '{32'h324db053};
/*############ DEBUG ############
test_input[30896:30903] = '{-59.2045278514, 66.4544526944, 4.38142004052, -49.5546348427, -57.9615493757, 85.2277988752, 66.1028168169, -24.3782805594};
test_label[3862] = '{85.2277988752};
test_output[3862] = '{1.19726620446e-08};
############ END DEBUG ############*/
test_input[30904:30911] = '{32'h41cedee3, 32'h42bb96cc, 32'h42814da7, 32'h414d9f8e, 32'h401c699d, 32'h42bfdfee, 32'h3e956fbb, 32'hc002d2e0};
test_label[3863] = '{32'h414d9f8e};
test_output[3863] = '{32'h42a664c8};
/*############ DEBUG ############
test_input[30904:30911] = '{25.8588319908, 93.7945235074, 64.6516652098, 12.8514535906, 2.4439460632, 95.9373610771, 0.291868054228, -2.04412076405};
test_label[3863] = '{12.8514535906};
test_output[3863] = '{83.1968417561};
############ END DEBUG ############*/
test_input[30912:30919] = '{32'h42a7d145, 32'hc1b0b55a, 32'hc298caab, 32'h3f3315cf, 32'h42a53207, 32'hc25de6a1, 32'hc200d00c, 32'h4183583e};
test_label[3864] = '{32'hc298caab};
test_output[3864] = '{32'h43208b11};
/*############ DEBUG ############
test_input[30912:30919] = '{83.9087309841, -22.0885499809, -76.3958380376, 0.699551495475, 82.5977069962, -55.4752252979, -32.2031703391, 16.4180860861};
test_label[3864] = '{-76.3958380376};
test_output[3864] = '{160.543226728};
############ END DEBUG ############*/
test_input[30920:30927] = '{32'hc24f2524, 32'h42add6e3, 32'h426e886f, 32'hc1bfa718, 32'hc05844ae, 32'hc20aae86, 32'h41dbe71a, 32'hc11305bb};
test_label[3865] = '{32'hc1bfa718};
test_output[3865] = '{32'h42ddc0a9};
/*############ DEBUG ############
test_input[30920:30927] = '{-51.7862712097, 86.91969739, 59.6332347725, -23.9565894, -3.37919176252, -34.6704316863, 27.4878419712, -9.18889863};
test_label[3865] = '{-23.9565894};
test_output[3865] = '{110.87628679};
############ END DEBUG ############*/
test_input[30928:30935] = '{32'hc0fb25aa, 32'hc20da680, 32'h42c10091, 32'h4270d708, 32'hc271e898, 32'hc2b04aa8, 32'h417c2acb, 32'hc2945434};
test_label[3866] = '{32'hc20da680};
test_output[3866] = '{32'h4303e9e9};
/*############ DEBUG ############
test_input[30928:30935] = '{-7.84834781273, -35.4125979631, 96.5011095653, 60.2099904311, -60.4771440372, -88.1458110342, 15.7604470462, -74.1644578146};
test_label[3866] = '{-35.4125979631};
test_output[3866] = '{131.913707528};
############ END DEBUG ############*/
test_input[30936:30943] = '{32'h429da37d, 32'h4297fbef, 32'h429c843b, 32'h42951d41, 32'hc1a2c5f2, 32'h426f8c8a, 32'hc0c0f08e, 32'h41f6be0a};
test_label[3867] = '{32'h429da37d};
test_output[3867] = '{32'h3efe7e26};
/*############ DEBUG ############
test_input[30936:30943] = '{78.8193120263, 75.9920554684, 78.258259671, 74.5571378446, -20.3466527111, 59.8872466229, -6.02936438591, 30.8427922638};
test_label[3867] = '{78.8193120263};
test_output[3867] = '{0.497056184706};
############ END DEBUG ############*/
test_input[30944:30951] = '{32'hc2a80b31, 32'h4279af3b, 32'hc28597aa, 32'h4280f888, 32'hc1c7b2c8, 32'hc1c255ff, 32'h42318191, 32'hc2500372};
test_label[3868] = '{32'h42318191};
test_output[3868] = '{32'h41a1d3b0};
/*############ DEBUG ############
test_input[30944:30951] = '{-84.0218614914, 62.4211228087, -66.7962200647, 64.4854127514, -24.9622953707, -24.291990747, 44.3765285837, -52.0033634624};
test_label[3868] = '{44.3765285837};
test_output[3868] = '{20.2283620975};
############ END DEBUG ############*/
test_input[30952:30959] = '{32'hc2bd8ba2, 32'h4284303f, 32'h42b12e25, 32'hc290d6b8, 32'hc104b866, 32'hc22f815f, 32'hc2005b8f, 32'h42830212};
test_label[3869] = '{32'hc2005b8f};
test_output[3869] = '{32'h42f15bec};
/*############ DEBUG ############
test_input[30952:30959] = '{-94.7727206296, 66.0942320467, 88.5901257887, -72.4193723584, -8.29501955363, -43.8763388708, -32.0894123833, 65.5040435692};
test_label[3869] = '{-32.0894123833};
test_output[3869] = '{120.679538172};
############ END DEBUG ############*/
test_input[30960:30967] = '{32'h41f102f2, 32'h423ff9ab, 32'h42213bcb, 32'h421cd30b, 32'h427b9085, 32'hc1d2c0d6, 32'h42a237db, 32'h42c6d1aa};
test_label[3870] = '{32'h42213bcb};
test_output[3870] = '{32'h426c6789};
/*############ DEBUG ############
test_input[30960:30967] = '{30.126438601, 47.9938160523, 40.3083914762, 39.2060959244, 62.8911339572, -26.3441572904, 81.1090951448, 99.4095016092};
test_label[3870] = '{40.3083914762};
test_output[3870] = '{59.1011101443};
############ END DEBUG ############*/
test_input[30968:30975] = '{32'hc19d2968, 32'hc2b1fa8c, 32'hc28e6372, 32'hc0133a3e, 32'h42b9bef6, 32'hc20be289, 32'hc23d27ae, 32'h41a66169};
test_label[3871] = '{32'hc2b1fa8c};
test_output[3871] = '{32'h4335dcc1};
/*############ DEBUG ############
test_input[30968:30975] = '{-19.6452180013, -88.989346422, -71.1942326399, -2.30042988809, 92.8729720011, -34.9712271903, -47.2887503786, 20.797562953};
test_label[3871] = '{-88.989346422};
test_output[3871] = '{181.862318423};
############ END DEBUG ############*/
test_input[30976:30983] = '{32'h42160667, 32'h4155b2e7, 32'hc0a8fc78, 32'h41bae129, 32'hc2aa94fa, 32'h3f630b31, 32'hc28f4a68, 32'h4149c718};
test_label[3872] = '{32'h42160667};
test_output[3872] = '{32'h3540d7be};
/*############ DEBUG ############
test_input[30976:30983] = '{37.5062537769, 13.3561775147, -5.2808189107, 23.3599414554, -85.2909725063, 0.886889493894, -71.6453274483, 12.6111071625};
test_label[3872] = '{37.5062537769};
test_output[3872] = '{7.18395213236e-07};
############ END DEBUG ############*/
test_input[30984:30991] = '{32'h41f5087d, 32'hc221d6cb, 32'h42190437, 32'h42c3618e, 32'hc1c671d8, 32'hc0d80025, 32'h413aee53, 32'hc289e046};
test_label[3873] = '{32'hc0d80025};
test_output[3873] = '{32'h42d0e190};
/*############ DEBUG ############
test_input[30984:30991] = '{30.6291439069, -40.4597598488, 38.254116806, 97.6905367874, -24.805587841, -6.75001759005, 11.6831847259, -68.9380337395};
test_label[3873] = '{-6.75001759005};
test_output[3873] = '{104.440554377};
############ END DEBUG ############*/
test_input[30992:30999] = '{32'hc1bbfc74, 32'h42bc9fcc, 32'h42a5699c, 32'h429625ce, 32'hc17b956b, 32'h42add51a, 32'hc299b9a3, 32'h428b4d51};
test_label[3874] = '{32'hc1bbfc74};
test_output[3874] = '{32'h42eb9f3a};
/*############ DEBUG ############
test_input[30992:30999] = '{-23.4982671916, 94.3120995936, 82.7062654961, 75.0738389731, -15.7239791371, 86.9162102965, -76.8625735597, 69.6510116805};
test_label[3874] = '{-23.4982671916};
test_output[3874] = '{117.810989479};
############ END DEBUG ############*/
test_input[31000:31007] = '{32'hc22f715f, 32'hc0f2e4ab, 32'hc0033bbe, 32'hc16ea818, 32'hc290e877, 32'h41fbc189, 32'h4284b0c5, 32'hc2999549};
test_label[3875] = '{32'hc290e877};
test_output[3875] = '{32'h430acc9e};
/*############ DEBUG ############
test_input[31000:31007] = '{-43.8607138944, -7.59041380004, -2.05052143261, -14.9160381359, -72.4540337097, 31.4694992991, 66.3452521296, -76.7915745094};
test_label[3875] = '{-72.4540337097};
test_output[3875] = '{138.799285839};
############ END DEBUG ############*/
test_input[31008:31015] = '{32'h3f557a66, 32'h4218d6de, 32'h42acdfac, 32'hc2a62e67, 32'hc243e5cb, 32'h42237c5f, 32'hc28ba10b, 32'h424840aa};
test_label[3876] = '{32'h42acdfac};
test_output[3876] = '{32'h25000000};
/*############ DEBUG ############
test_input[31008:31015] = '{0.833898908291, 38.2098317745, 86.4368561726, -83.0906320827, -48.9744056597, 40.8714556978, -69.81453679, 50.0631475835};
test_label[3876] = '{86.4368561726};
test_output[3876] = '{1.11022302463e-16};
############ END DEBUG ############*/
test_input[31016:31023] = '{32'hc2b4fe9d, 32'h41a5fe97, 32'h41cc0d52, 32'hc2b19ba2, 32'hc2052b0d, 32'hc071f5df, 32'hc29b23b5, 32'hc24cb31b};
test_label[3877] = '{32'h41a5fe97};
test_output[3877] = '{32'h40988100};
/*############ DEBUG ############
test_input[31016:31023] = '{-90.4972925679, 20.7493107467, 25.5065048758, -88.8039679152, -33.2920412148, -3.78063185487, -77.5697404814, -51.1749076848};
test_label[3877] = '{20.7493107467};
test_output[3877] = '{4.76574712481};
############ END DEBUG ############*/
test_input[31024:31031] = '{32'hc1c22c61, 32'hc2bbbdb9, 32'hc2976a59, 32'hc23ef811, 32'h427fdbe9, 32'h4293e428, 32'hc21c7d71, 32'h4286732e};
test_label[3878] = '{32'h4286732e};
test_output[3878] = '{32'h40d719d9};
/*############ DEBUG ############
test_input[31024:31031] = '{-24.271669127, -93.8705491628, -75.7077071351, -47.7422528934, 63.964756795, 73.9456153291, -39.122499859, 67.2249611827};
test_label[3878] = '{67.2249611827};
test_output[3878] = '{6.72190538987};
############ END DEBUG ############*/
test_input[31032:31039] = '{32'h40f199c5, 32'hc1c39be2, 32'hc1b868fa, 32'hc23d4dd5, 32'h429f7f2c, 32'hc2bedd5f, 32'h42939fc4, 32'hc2a69886};
test_label[3879] = '{32'hc1c39be2};
test_output[3879] = '{32'h42d0677e};
/*############ DEBUG ############
test_input[31032:31039] = '{7.55002065331, -24.4511153536, -23.0512586301, -47.3260085644, 79.7483804974, -95.4323638961, 73.8120443203, -83.2978975033};
test_label[3879] = '{-24.4511153536};
test_output[3879] = '{104.202134059};
############ END DEBUG ############*/
test_input[31040:31047] = '{32'h4299c855, 32'h4296ded9, 32'h423eed4e, 32'h428f2a5f, 32'hc2c1a04c, 32'hc2aa7219, 32'h42c692ae, 32'h42b60f6d};
test_label[3880] = '{32'h423eed4e};
test_output[3880] = '{32'h424e3852};
/*############ DEBUG ############
test_input[31040:31047] = '{76.8912760672, 75.4352489017, 47.7317416449, 71.5827526913, -96.8130807552, -85.2228491815, 99.2864815214, 91.0301265058};
test_label[3880] = '{47.7317416449};
test_output[3880] = '{51.5549994466};
############ END DEBUG ############*/
test_input[31048:31055] = '{32'h40cce12d, 32'hc26a8c38, 32'h42454ff8, 32'hc2c4d245, 32'hc2a9c23d, 32'h40e1e612, 32'h42293687, 32'h4219f56d};
test_label[3881] = '{32'h40cce12d};
test_output[3881] = '{32'h422bb4c1};
/*############ DEBUG ############
test_input[31048:31055] = '{6.40248741324, -58.6369332153, 49.3280955736, -98.4106828425, -84.879370448, 7.05933493151, 42.3032505116, 38.489673374};
test_label[3881] = '{6.40248741324};
test_output[3881] = '{42.9265168832};
############ END DEBUG ############*/
test_input[31056:31063] = '{32'hc28f51f7, 32'hc251e906, 32'h426944a0, 32'hc2361fcb, 32'hc267ffa8, 32'hc157a2c8, 32'hc1c6d72c, 32'h414cb591};
test_label[3882] = '{32'hc1c6d72c};
test_output[3882] = '{32'h42a6581b};
/*############ DEBUG ############
test_input[31056:31063] = '{-71.6600903386, -52.4775617978, 58.3170178749, -45.531048492, -57.9996651049, -13.4772411855, -24.8550640136, 12.7943278984};
test_label[3882] = '{-24.8550640136};
test_output[3882] = '{83.1720818885};
############ END DEBUG ############*/
test_input[31064:31071] = '{32'h4212d284, 32'hc1a84032, 32'hc24b3324, 32'h424c8ded, 32'h42128616, 32'h42b5d493, 32'hc2202abe, 32'h411d4f94};
test_label[3883] = '{32'h42b5d493};
test_output[3883] = '{32'h80000000};
/*############ DEBUG ############
test_input[31064:31071] = '{36.7055835526, -21.0313445128, -50.7999405925, 51.1385986905, 36.630942164, 90.915183198, -40.0417390075, 9.83192872707};
test_label[3883] = '{90.915183198};
test_output[3883] = '{-0.0};
############ END DEBUG ############*/
test_input[31072:31079] = '{32'hc2b1d8b2, 32'hc17380bf, 32'hc288c118, 32'hbf3e404b, 32'h4280b957, 32'h40b2fa5f, 32'h42a66e6b, 32'hc09be270};
test_label[3884] = '{32'hc09be270};
test_output[3884] = '{32'h42b02c92};
/*############ DEBUG ############
test_input[31072:31079] = '{-88.9232363759, -15.218932566, -68.3771326349, -0.743168548643, 64.3619944849, 5.59306301525, 83.2156590035, -4.87139121596};
test_label[3884] = '{-4.87139121596};
test_output[3884] = '{88.0870502259};
############ END DEBUG ############*/
test_input[31080:31087] = '{32'hc26b89b5, 32'h41a7a6b8, 32'h428224f8, 32'h422405c3, 32'h42b0d1a7, 32'hc2185373, 32'h42c05266, 32'h41742076};
test_label[3885] = '{32'hc2185373};
test_output[3885] = '{32'h43063e2c};
/*############ DEBUG ############
test_input[31080:31087] = '{-58.8844810085, 20.9564062084, 65.0722070388, 41.005628463, 88.4094771809, -38.0814925263, 96.1609369188, 15.2579253376};
test_label[3885] = '{-38.0814925263};
test_output[3885] = '{134.242859467};
############ END DEBUG ############*/
test_input[31088:31095] = '{32'hc272c3dd, 32'hc24101c4, 32'hc29cc0eb, 32'hc1c11f5b, 32'hc1b8e60c, 32'hc291ef27, 32'h423bae6f, 32'h4045e750};
test_label[3886] = '{32'h423bae6f};
test_output[3886] = '{32'h80000000};
/*############ DEBUG ############
test_input[31088:31095] = '{-60.6912724705, -48.2517243142, -78.3767893291, -24.140311188, -23.1123272667, -72.9670963469, 46.9203456675, 3.09224316896};
test_label[3886] = '{46.9203456675};
test_output[3886] = '{-0.0};
############ END DEBUG ############*/
test_input[31096:31103] = '{32'h428b8cc5, 32'h42472442, 32'hc1e8f7d2, 32'hc2c7ffdc, 32'hc223900f, 32'hc27f0d0a, 32'hc1bf3c58, 32'hc032762b};
test_label[3887] = '{32'hc27f0d0a};
test_output[3887] = '{32'h430589a5};
/*############ DEBUG ############
test_input[31096:31103] = '{69.7749392573, 49.7854089864, -29.1210065724, -99.9997291488, -40.8906829823, -63.7627338074, -23.9044654812, -2.78846228806};
test_label[3887] = '{-63.7627338074};
test_output[3887] = '{133.537673067};
############ END DEBUG ############*/
test_input[31104:31111] = '{32'hc2bda7a2, 32'h3f4f48ff, 32'h42038f8d, 32'hc24b473b, 32'h428a1e55, 32'hc2823a27, 32'h409204c7, 32'h40ed7dea};
test_label[3888] = '{32'hc2823a27};
test_output[3888] = '{32'h43062c3e};
/*############ DEBUG ############
test_input[31104:31111] = '{-94.8274113547, 0.809707598004, 32.8901866098, -50.8195591066, 69.0592393529, -65.1135812823, 4.56308317744, 7.42162048545};
test_label[3888] = '{-65.1135812823};
test_output[3888] = '{134.172820635};
############ END DEBUG ############*/
test_input[31112:31119] = '{32'hc29def65, 32'hc215a3d1, 32'h428d7857, 32'h42c43d3a, 32'hc219be7e, 32'h423c41ae, 32'h41f995f8, 32'h4089260c};
test_label[3889] = '{32'hc219be7e};
test_output[3889] = '{32'h43088e3c};
/*############ DEBUG ############
test_input[31112:31119] = '{-78.9675711842, -37.4099763076, 70.7350413524, 98.1195815847, -38.4360272463, 47.0641390886, 31.1982274569, 4.28589456942};
test_label[3889] = '{-38.4360272463};
test_output[3889] = '{136.555608831};
############ END DEBUG ############*/
test_input[31120:31127] = '{32'hc29e382e, 32'hc20966cd, 32'h4271584e, 32'hc1feac9d, 32'h424fd9ca, 32'h405d921b, 32'h42940d79, 32'h42c3e3b0};
test_label[3890] = '{32'hc29e382e};
test_output[3890] = '{32'h43310def};
/*############ DEBUG ############
test_input[31120:31127] = '{-79.1097285612, -34.3503908927, 60.3362355854, -31.8342843947, 51.962686095, 3.46204253156, 74.0263153755, 97.9447057289};
test_label[3890] = '{-79.1097285612};
test_output[3890] = '{177.05443429};
############ END DEBUG ############*/
test_input[31128:31135] = '{32'h41aaf1d0, 32'hc1d2fd2c, 32'h42c0637b, 32'h428e4a06, 32'h426adfd2, 32'h4298f500, 32'h42afa1e9, 32'h424f95a2};
test_label[3891] = '{32'h4298f500};
test_output[3891] = '{32'h419dba64};
/*############ DEBUG ############
test_input[31128:31135] = '{21.3680719417, -26.3736198812, 96.194295349, 71.1445759878, 58.7185760169, 76.4785148627, 87.8162316984, 51.8961245381};
test_label[3891] = '{76.4785148627};
test_output[3891] = '{19.7160103172};
############ END DEBUG ############*/
test_input[31136:31143] = '{32'h4213f7ce, 32'hc2597f46, 32'h42c7f2ac, 32'hc2b5e8bb, 32'hc129291d, 32'hc243253d, 32'hc251760e, 32'hc2969e48};
test_label[3892] = '{32'h4213f7ce};
test_output[3892] = '{32'h427bed89};
/*############ DEBUG ############
test_input[31136:31143] = '{36.9919981505, -54.3742907834, 99.9739661505, -90.9545482001, -10.5725378771, -48.7863673169, -52.3652881493, -75.309144571};
test_label[3892] = '{36.9919981505};
test_output[3892] = '{62.981968};
############ END DEBUG ############*/
test_input[31144:31151] = '{32'hc1a84477, 32'h419076fa, 32'hc1737ae6, 32'h425e49c1, 32'hc28306ad, 32'hc20779a9, 32'h40db37c6, 32'hc20f8755};
test_label[3893] = '{32'h425e49c1};
test_output[3893] = '{32'h80000000};
/*############ DEBUG ############
test_input[31144:31151] = '{-21.0334296114, 18.0580935478, -15.2175045176, 55.5720265097, -65.5130406722, -33.8688103451, 6.85055836193, -35.8821616477};
test_label[3893] = '{55.5720265097};
test_output[3893] = '{-0.0};
############ END DEBUG ############*/
test_input[31152:31159] = '{32'hc1e39099, 32'hc29ff516, 32'h4176f027, 32'h42b64ac5, 32'h428904c5, 32'hc2b6fa90, 32'hc2c470f4, 32'hc23a523a};
test_label[3894] = '{32'h4176f027};
test_output[3894] = '{32'h42976cc0};
/*############ DEBUG ############
test_input[31152:31159] = '{-28.4456036131, -79.9786865687, 15.4336309255, 91.1460357994, 68.5093161437, -91.4893796598, -98.2206122149, -46.5802998473};
test_label[3894] = '{15.4336309255};
test_output[3894] = '{75.712404874};
############ END DEBUG ############*/
test_input[31160:31167] = '{32'h42bb0b64, 32'hc0adf10f, 32'hc064f56f, 32'h4295e902, 32'hc22ef1ad, 32'hc21062fd, 32'hc2666963, 32'hc2a0cb63};
test_label[3895] = '{32'hc22ef1ad};
test_output[3895] = '{32'h4309421d};
/*############ DEBUG ############
test_input[31160:31167] = '{93.5222453528, -5.4356761576, -3.57747999109, 74.9550900663, -43.7360104706, -36.0966683963, -57.6029164397, -80.3972427971};
test_label[3895] = '{-43.7360104706};
test_output[3895] = '{137.258255832};
############ END DEBUG ############*/
test_input[31168:31175] = '{32'hc26aa0f9, 32'hc290d3e0, 32'hc276ce9a, 32'hc250cf0c, 32'h42c0acc4, 32'h42c4d807, 32'h41b22858, 32'hc1d14fa4};
test_label[3896] = '{32'hc290d3e0};
test_output[3896] = '{32'h432af3f6};
/*############ DEBUG ############
test_input[31168:31175] = '{-58.6571985346, -72.4138203169, -61.7017591647, -52.2021946367, 96.3374306404, 98.4219314803, 22.2696988241, -26.1638878324};
test_label[3896] = '{-72.4138203169};
test_output[3896] = '{170.952973951};
############ END DEBUG ############*/
test_input[31176:31183] = '{32'hc237c856, 32'hc2b6ffd6, 32'h3f5e7e78, 32'hc13d96a9, 32'hc2c79e22, 32'hc1ac176e, 32'hc1774e38, 32'hc2c0498e};
test_label[3897] = '{32'hc13d96a9};
test_output[3897] = '{32'h414b7e94};
/*############ DEBUG ############
test_input[31176:31183] = '{-45.9456397813, -91.4996797385, 0.869117254849, -11.8492822749, -99.8088565573, -21.5114400774, -15.4565961664, -96.1436630766};
test_label[3897] = '{-11.8492822749};
test_output[3897] = '{12.7184026067};
############ END DEBUG ############*/
test_input[31184:31191] = '{32'h4163c63e, 32'hc2155ea1, 32'h4239d88a, 32'h41b60252, 32'h41210542, 32'h42a8cf42, 32'hc26a07e3, 32'h41f88272};
test_label[3898] = '{32'h4239d88a};
test_output[3898] = '{32'h4217c5fa};
/*############ DEBUG ############
test_input[31184:31191] = '{14.2358990501, -37.342410497, 46.4614647172, 22.7511326485, 10.0637833971, 84.4047997092, -58.5077019467, 31.0636939311};
test_label[3898] = '{46.4614647172};
test_output[3898] = '{37.943334992};
############ END DEBUG ############*/
test_input[31192:31199] = '{32'hc2558704, 32'hc18f19f9, 32'h418d2e02, 32'hc21d35d2, 32'hc1b39fa2, 32'hc284d05a, 32'hc05b47a2, 32'h428f77c6};
test_label[3899] = '{32'hc1b39fa2};
test_output[3899] = '{32'h42bc5faf};
/*############ DEBUG ############
test_input[31192:31199] = '{-53.3818511524, -17.8876822622, 17.6474647628, -39.3025580163, -22.452945457, -66.4069347144, -3.4262470385, 71.7339340226};
test_label[3899] = '{-22.452945457};
test_output[3899] = '{94.1868794796};
############ END DEBUG ############*/
test_input[31200:31207] = '{32'h42860779, 32'hc2844c3b, 32'h4235365e, 32'h4252d571, 32'h41d9223e, 32'hc231f808, 32'h42c28e0b, 32'hc2282f2c};
test_label[3900] = '{32'h41d9223e};
test_output[3900] = '{32'h428c457b};
/*############ DEBUG ############
test_input[31200:31207] = '{67.0145977152, -66.1488844367, 45.3030938262, 52.7084403045, 27.1417198927, -44.4922165657, 97.2774264638, -42.0460648671};
test_label[3900] = '{27.1417198927};
test_output[3900] = '{70.135706571};
############ END DEBUG ############*/
test_input[31208:31215] = '{32'hc20b5abe, 32'h422a1096, 32'hc1860647, 32'hc2b34e70, 32'hc28317a5, 32'hc20cda59, 32'hc2a9e713, 32'h41e8751a};
test_label[3901] = '{32'h41e8751a};
test_output[3901] = '{32'h41575823};
/*############ DEBUG ############
test_input[31208:31215] = '{-34.8386154801, 42.5161954048, -16.7530655346, -89.6531945862, -65.5461789219, -35.2132309874, -84.9513152246, 29.0571788879};
test_label[3901] = '{29.0571788879};
test_output[3901] = '{13.4590179451};
############ END DEBUG ############*/
test_input[31216:31223] = '{32'h40e2e020, 32'hc260e321, 32'h41d2115b, 32'h42516edc, 32'h424e1392, 32'h4285cef8, 32'h4198d31b, 32'h41e1b650};
test_label[3902] = '{32'hc260e321};
test_output[3902] = '{32'h42f64089};
/*############ DEBUG ############
test_input[31216:31223] = '{7.08985899382, -56.2218046195, 26.2584734304, 52.3582601111, 51.5191127699, 66.9042386209, 19.1030797408, 28.2140202128};
test_label[3902] = '{-56.2218046195};
test_output[3902] = '{123.12604393};
############ END DEBUG ############*/
test_input[31224:31231] = '{32'h41a0e438, 32'hc2bd62a4, 32'h41d98617, 32'h41d47a6a, 32'hc2a8c4db, 32'h42b6c59b, 32'hc26426ac, 32'hc10f9062};
test_label[3903] = '{32'hc2bd62a4};
test_output[3903] = '{32'h433a141f};
/*############ DEBUG ############
test_input[31224:31231] = '{20.1114342226, -94.6926587135, 27.1904739372, 26.5597719476, -84.3844868504, 91.3859462745, -57.0377643258, -8.97274995483};
test_label[3903] = '{-94.6926587135};
test_output[3903] = '{186.078604988};
############ END DEBUG ############*/
test_input[31232:31239] = '{32'h42bf66bf, 32'hc22e6b34, 32'h4274e4ec, 32'hc2815737, 32'hc0d75590, 32'h4239be76, 32'h420be6f0, 32'hc1107d82};
test_label[3904] = '{32'hc22e6b34};
test_output[3904] = '{32'h430b4e2d};
/*############ DEBUG ############
test_input[31232:31239] = '{95.7006771288, -43.6046898147, 61.2235561786, -64.6703393531, -6.72919462874, 46.4359973204, 34.9755233195, -9.03064201293};
test_label[3904] = '{-43.6046898147};
test_output[3904] = '{139.305366944};
############ END DEBUG ############*/
test_input[31240:31247] = '{32'hc2bfc96d, 32'h424ae2dd, 32'h40482c8a, 32'h42a08866, 32'hc2813d5b, 32'hc2813035, 32'h42b174ec, 32'h41dd369b};
test_label[3905] = '{32'hc2813035};
test_output[3905] = '{32'h4319529e};
/*############ DEBUG ############
test_input[31240:31247] = '{-95.8934086072, 50.7215479074, 3.12771847245, 80.2664042424, -64.6198354203, -64.5941553375, 88.7283599435, 27.6516627811};
test_label[3905] = '{-64.5941553375};
test_output[3905] = '{153.322726617};
############ END DEBUG ############*/
test_input[31248:31255] = '{32'h42a73936, 32'h4262dd33, 32'hc1a6a369, 32'h4284118a, 32'h3f96dd1c, 32'h4220eb72, 32'h40d42359, 32'h3fa9a31e};
test_label[3906] = '{32'h4220eb72};
test_output[3906] = '{32'h422d86fa};
/*############ DEBUG ############
test_input[31248:31255] = '{83.6117396818, 56.7160135267, -20.8297909759, 66.034257425, 1.17862277331, 40.2299274264, 6.62931502764, 1.3252904423};
test_label[3906] = '{40.2299274264};
test_output[3906] = '{43.3818122786};
############ END DEBUG ############*/
test_input[31256:31263] = '{32'hc28373ab, 32'hc29e886f, 32'h4248263f, 32'h428ce716, 32'hc24c3018, 32'h406c11b5, 32'h4241f928, 32'h42a80dfa};
test_label[3907] = '{32'hc29e886f};
test_output[3907] = '{32'h43234b34};
/*############ DEBUG ############
test_input[31256:31263] = '{-65.7259176665, -79.2664683444, 50.0373491974, 70.4513371371, -51.0469664791, 3.68858063344, 48.4933164631, 84.0272958659};
test_label[3907] = '{-79.2664683444};
test_output[3907] = '{163.293765481};
############ END DEBUG ############*/
test_input[31264:31271] = '{32'hc05313c8, 32'h426696c5, 32'hc1419a87, 32'h42376aee, 32'hc2751c00, 32'hc19fdd8f, 32'hc22a0bd4, 32'hc288a69a};
test_label[3908] = '{32'hc19fdd8f};
test_output[3908] = '{32'h429b42c7};
/*############ DEBUG ############
test_input[31264:31271] = '{-3.2980824081, 57.6472361253, -12.1002260204, 45.8544247556, -61.2773437355, -19.983182607, -42.5115509622, -68.3253926817};
test_label[3908] = '{-19.983182607};
test_output[3908] = '{77.630426291};
############ END DEBUG ############*/
test_input[31272:31279] = '{32'h41bd9cbf, 32'h42838497, 32'h4297ccf8, 32'h42220984, 32'hc223cfc5, 32'hc23559c6, 32'hc23aa985, 32'hc29c35c4};
test_label[3909] = '{32'hc29c35c4};
test_output[3909] = '{32'h431a0160};
/*############ DEBUG ############
test_input[31272:31279] = '{23.7015353891, 65.7589608731, 75.9003274194, 40.5092944778, -40.9529001417, -45.3376678853, -46.6655460468, -78.1050071761};
test_label[3909] = '{-78.1050071761};
test_output[3909] = '{154.00537401};
############ END DEBUG ############*/
test_input[31280:31287] = '{32'hc274deb6, 32'hc215d802, 32'hc2878df1, 32'h42829460, 32'h3dba8963, 32'hc29e2a59, 32'hc1d2dbee, 32'h42657cf4};
test_label[3910] = '{32'hc29e2a59};
test_output[3910] = '{32'h43105f74};
/*############ DEBUG ############
test_input[31280:31287] = '{-61.2174912839, -37.4609463122, -67.7772314584, 65.2897936319, 0.0910823579603, -79.0827130124, -26.3573873255, 57.3720230504};
test_label[3910] = '{-79.0827130124};
test_output[3910] = '{144.372870791};
############ END DEBUG ############*/
test_input[31288:31295] = '{32'hc29a4487, 32'hc2bb8e2d, 32'hc2bc2729, 32'h409707d7, 32'h425dd620, 32'hc2a65f2f, 32'h42a5cb6e, 32'h4233b746};
test_label[3911] = '{32'h4233b746};
test_output[3911] = '{32'h4217df96};
/*############ DEBUG ############
test_input[31288:31295] = '{-77.1338459787, -93.7776858793, -94.0764811077, 4.71970712447, 55.459104833, -83.1859018542, 82.8973239592, 44.9289773315};
test_label[3911] = '{44.9289773315};
test_output[3911] = '{37.9683466278};
############ END DEBUG ############*/
test_input[31296:31303] = '{32'hc2a2a884, 32'hc2b57730, 32'hc2aa5c59, 32'h42b2316f, 32'h41548cae, 32'hc2725db5, 32'h426a6f6d, 32'h42ad9e54};
test_label[3912] = '{32'hc2725db5};
test_output[3912] = '{32'h4315c8e7};
/*############ DEBUG ############
test_input[31296:31303] = '{-81.3291335297, -90.7327847704, -85.1803680448, 89.0965513263, 13.2843456767, -60.5915116277, 58.6088145826, 86.8092331934};
test_label[3912] = '{-60.5915116277};
test_output[3912] = '{149.784770711};
############ END DEBUG ############*/
test_input[31304:31311] = '{32'hc29f1aab, 32'hc2ab48cd, 32'hc1379fd4, 32'h42509003, 32'hc20d7ec4, 32'h42aefe64, 32'h41952bf6, 32'hc28bbdb1};
test_label[3913] = '{32'h42509003};
test_output[3913] = '{32'h420d6cc6};
/*############ DEBUG ############
test_input[31304:31311] = '{-79.5520852664, -85.6421886373, -11.4765203331, 52.14063713, -35.3737947958, 87.4968598755, 18.6464643939, -69.8704943652};
test_label[3913] = '{52.14063713};
test_output[3913] = '{35.3562227455};
############ END DEBUG ############*/
test_input[31312:31319] = '{32'hc186248b, 32'h421c65a8, 32'h41ccf454, 32'hc2b0ad44, 32'hc255cb0e, 32'hc20f6811, 32'h42baac60, 32'h412ffbfc};
test_label[3914] = '{32'hc255cb0e};
test_output[3914] = '{32'h4312c8f4};
/*############ DEBUG ############
test_input[31312:31319] = '{-16.7678428325, 39.0992743566, 25.6193003689, -88.3384057846, -53.4482946789, -35.8516268085, 93.336673194, 10.9990198144};
test_label[3914] = '{-53.4482946789};
test_output[3914] = '{146.784967873};
############ END DEBUG ############*/
test_input[31320:31327] = '{32'h422657e5, 32'h4286a291, 32'hc1ab7870, 32'h42999ac9, 32'hc22377c9, 32'hc2b20cb7, 32'hc18ab05a, 32'hc16b4158};
test_label[3915] = '{32'hc22377c9};
test_output[3915] = '{32'h42eb56b8};
/*############ DEBUG ############
test_input[31320:31327] = '{41.5858361464, 67.3175106033, -21.4338076033, 76.8023183267, -40.8669773336, -89.0248314762, -17.3361100832, -14.7034534403};
test_label[3915] = '{-40.8669773336};
test_output[3915] = '{117.669371655};
############ END DEBUG ############*/
test_input[31328:31335] = '{32'hc2af69f4, 32'hc23fceb7, 32'hc2931acf, 32'h421f8689, 32'h42059068, 32'h41862085, 32'h425e1fd8, 32'hc2a8b3c4};
test_label[3916] = '{32'h425e1fd8};
test_output[3916] = '{32'h342bc7c0};
/*############ DEBUG ############
test_input[31328:31335] = '{-87.7069404911, -47.9518698438, -73.5523636383, 39.8813824662, 33.3910198391, 16.7658796049, 55.531098455, -84.3511057753};
test_label[3916] = '{55.531098455};
test_output[3916] = '{1.59982848998e-07};
############ END DEBUG ############*/
test_input[31336:31343] = '{32'hc249716c, 32'hc037b274, 32'hc2c33286, 32'hc22aad4c, 32'hc255f583, 32'h404890e5, 32'h40f2d5d4, 32'hc2978082};
test_label[3917] = '{32'hc22aad4c};
test_output[3917] = '{32'h424913e3};
/*############ DEBUG ############
test_input[31336:31343] = '{-50.3607642556, -2.87026690661, -97.5986818709, -42.6692354723, -53.4897563963, 3.13384370103, 7.58860201868, -75.7509909857};
test_label[3917] = '{-42.6692354723};
test_output[3917] = '{50.2694219526};
############ END DEBUG ############*/
test_input[31344:31351] = '{32'hbec2307c, 32'h429d2ecb, 32'hc2b38764, 32'hc24073e8, 32'h42963d44, 32'hc2a5f114, 32'h41f4d597, 32'h42ad7dc3};
test_label[3918] = '{32'hc2b38764};
test_output[3918] = '{32'h433082a7};
/*############ DEBUG ############
test_input[31344:31351] = '{-0.379276169812, 78.5913960541, -89.7644368399, -48.1131885647, 75.1196584778, -82.9708555116, 30.6042925435, 86.7456263845};
test_label[3918] = '{-89.7644368399};
test_output[3918] = '{176.510359628};
############ END DEBUG ############*/
test_input[31352:31359] = '{32'h428444ea, 32'hc28ab793, 32'hc21959d7, 32'h40bc1d26, 32'h3f39abd9, 32'hc2c3a065, 32'hc0ff0df5, 32'hbf274136};
test_label[3919] = '{32'hc2c3a065};
test_output[3919] = '{32'h4323f2a7};
/*############ DEBUG ############
test_input[31352:31359] = '{66.1345972064, -69.3585420685, -38.3377348352, 5.87855826845, 0.725278458348, -97.8132681816, -7.97045361912, -0.653338768422};
test_label[3919] = '{-97.8132681816};
test_output[3919] = '{163.947865388};
############ END DEBUG ############*/
test_input[31360:31367] = '{32'hc181db42, 32'hc2b78518, 32'h420486ef, 32'h4234b82c, 32'h42bf2151, 32'hc2935ebc, 32'hc11342c9, 32'hc168257c};
test_label[3920] = '{32'hc168257c};
test_output[3920] = '{32'h42dc2600};
/*############ DEBUG ############
test_input[31360:31367] = '{-16.232059525, -91.7599509789, 33.1317701372, 45.1798561715, 95.565068074, -73.6850248061, -9.20380542786, -14.509151455};
test_label[3920] = '{-14.509151455};
test_output[3920] = '{110.074219529};
############ END DEBUG ############*/
test_input[31368:31375] = '{32'hc2c2d77f, 32'h42b2af27, 32'h422aad5f, 32'h423e58df, 32'h429d99b1, 32'h41bd07c9, 32'hc22dc59e, 32'hc24ce1cd};
test_label[3921] = '{32'h42b2af27};
test_output[3921] = '{32'h37dd81c1};
/*############ DEBUG ############
test_input[31368:31375] = '{-97.4208899796, 89.3420965361, 42.669307388, 47.5867896436, 78.8001781101, 23.6288010675, -43.4429849684, -51.2205068925};
test_label[3921] = '{89.3420965361};
test_output[3921] = '{2.64056744708e-05};
############ END DEBUG ############*/
test_input[31376:31383] = '{32'h418e9fcf, 32'hc19879da, 32'h4287ef87, 32'hc269cea7, 32'hc1096ef5, 32'hc29c68e1, 32'hc1ca5024, 32'h42ab44e3};
test_label[3922] = '{32'hc269cea7};
test_output[3922] = '{32'h4310161b};
/*############ DEBUG ############
test_input[31376:31383] = '{17.8280315468, -19.0594981188, 67.9678243828, -58.4518095857, -8.58958903473, -78.2048427286, -25.2891313861, 85.6345410484};
test_label[3922] = '{-58.4518095857};
test_output[3922] = '{144.086350655};
############ END DEBUG ############*/
test_input[31384:31391] = '{32'h42831f52, 32'h42b683af, 32'h422cbcec, 32'h41fce1bb, 32'h42452fb1, 32'hc2998cec, 32'hc29b9c8c, 32'hc21f05ca};
test_label[3923] = '{32'h42b683af};
test_output[3923] = '{32'h2cf39e00};
/*############ DEBUG ############
test_input[31384:31391] = '{65.5611697642, 91.257197673, 43.1844955775, 31.6102194434, 49.2965722631, -76.7752416463, -77.8057583912, -39.7556539507};
test_label[3923] = '{91.257197673};
test_output[3923] = '{6.9240169154e-12};
############ END DEBUG ############*/
test_input[31392:31399] = '{32'hc064fe63, 32'h410d0d0e, 32'h4206903b, 32'hc203c51a, 32'h424fb5e2, 32'hc2b596ed, 32'h410a3583, 32'hc2975a36};
test_label[3924] = '{32'hc203c51a};
test_output[3924] = '{32'h42a9bd7e};
/*############ DEBUG ############
test_input[31392:31399] = '{-3.57802654448, 8.81568697384, 33.6408513889, -32.9424827592, 51.9276185908, -90.7947768657, 8.63806400455, -75.6761922609};
test_label[3924] = '{-32.9424827592};
test_output[3924] = '{84.8701013614};
############ END DEBUG ############*/
test_input[31400:31407] = '{32'h4287c820, 32'h41d887c4, 32'h4294e66c, 32'h42193d1e, 32'h4281992d, 32'hc23b9883, 32'h4287794a, 32'hc1af716e};
test_label[3925] = '{32'h41d887c4};
test_output[3925] = '{32'h423d8bb7};
/*############ DEBUG ############
test_input[31400:31407] = '{67.8908653996, 27.0662921677, 74.4500404259, 38.309685021, 64.7991679395, -46.8989386624, 67.736889704, -21.9303853735};
test_label[3925] = '{27.0662921677};
test_output[3925] = '{47.3864408839};
############ END DEBUG ############*/
test_input[31408:31415] = '{32'h40e3bc35, 32'hc26275c2, 32'hc283c068, 32'hc11a703c, 32'hc28b7afc, 32'h42ab9708, 32'hc2ad2884, 32'h4253fbdc};
test_label[3926] = '{32'hc28b7afc};
test_output[3926] = '{32'h431b8902};
/*############ DEBUG ############
test_input[31408:31415] = '{7.11672456361, -56.6149978777, -65.8757906246, -9.65240129611, -69.7402001345, 85.7949833978, -86.5791328576, 52.9959582162};
test_label[3926] = '{-69.7402001345};
test_output[3926] = '{155.535183532};
############ END DEBUG ############*/
test_input[31416:31423] = '{32'hc293bda7, 32'hc1ce5ab0, 32'h4266fcd0, 32'hc2a18331, 32'hc2ab6d3f, 32'hc2a1989d, 32'h40d5ca27, 32'h4268dc44};
test_label[3927] = '{32'hc2a1989d};
test_output[3927] = '{32'h430b7fd7};
/*############ DEBUG ############
test_input[31416:31423] = '{-73.870412314, -25.7942817731, 57.7468856781, -80.7562341324, -85.7133706576, -80.7980736851, 6.68092656388, 58.2151034893};
test_label[3927] = '{-80.7980736851};
test_output[3927] = '{139.499372221};
############ END DEBUG ############*/
test_input[31424:31431] = '{32'h40862132, 32'hc1cedc1c, 32'h41aa0d60, 32'hc07ce10b, 32'h41c63d9d, 32'h4214159a, 32'h4262e5e1, 32'h41d1e236};
test_label[3928] = '{32'h41c63d9d};
test_output[3928] = '{32'h41ff8e26};
/*############ DEBUG ############
test_input[31424:31431] = '{4.19155234473, -25.8574745811, 21.2565300678, -3.95123543201, 24.7800836883, 37.0210967159, 56.7244929236, 26.2354541671};
test_label[3928] = '{24.7800836883};
test_output[3928] = '{31.9444092381};
############ END DEBUG ############*/
test_input[31432:31439] = '{32'hc294216b, 32'h42aee636, 32'h42139185, 32'h41b35b22, 32'h41c5528f, 32'h423f6327, 32'h42bda38c, 32'h418dd8ef};
test_label[3929] = '{32'h42aee636};
test_output[3929] = '{32'h40ebda86};
/*############ DEBUG ############
test_input[31432:31439] = '{-74.0652674723, 87.4496302059, 36.8921083041, 22.419498553, 24.6653126148, 47.8468285834, 94.8194258301, 17.7309250297};
test_label[3929] = '{87.4496302059};
test_output[3929] = '{7.3704254228};
############ END DEBUG ############*/
test_input[31440:31447] = '{32'h42bd4922, 32'h427a4e4b, 32'h42b7e673, 32'h424b7f02, 32'h42b3fc14, 32'hc21970f1, 32'h41a91445, 32'h427968a2};
test_label[3930] = '{32'h42b3fc14};
test_output[3930] = '{32'h40973277};
/*############ DEBUG ############
test_input[31440:31447] = '{94.6428388669, 62.5764569624, 91.9500991684, 50.8740295691, 89.9923422671, -38.3602939534, 21.1348969844, 62.3521798784};
test_label[3930] = '{89.9923422671};
test_output[3930] = '{4.72491002386};
############ END DEBUG ############*/
test_input[31448:31455] = '{32'h3ee2cbc1, 32'h413aa42f, 32'hbf3cd4bb, 32'hc2436806, 32'hc1811da9, 32'h4231f607, 32'hc29ae84b, 32'hc2b58359};
test_label[3931] = '{32'hbf3cd4bb};
test_output[3931] = '{32'h4234e95a};
/*############ DEBUG ############
test_input[31448:31455] = '{0.442960761499, 11.6650839919, -0.737621009127, -48.8515869878, -16.1394827409, 44.4902608384, -77.4536983243, -90.7565417345};
test_label[3931] = '{-0.737621009127};
test_output[3931] = '{45.2278818475};
############ END DEBUG ############*/
test_input[31456:31463] = '{32'h428e675d, 32'hc28a6988, 32'hc2b37e93, 32'h4242ddb0, 32'h4276c649, 32'h42ae3044, 32'hc18c164b, 32'hc25425da};
test_label[3932] = '{32'hc28a6988};
test_output[3932] = '{32'h431c4ce6};
/*############ DEBUG ############
test_input[31456:31463] = '{71.2018836658, -69.2061135582, -89.7472164929, 48.716490919, 61.6936373413, 87.09426973, -17.5108859188, -53.036963399};
test_label[3932] = '{-69.2061135582};
test_output[3932] = '{156.300383414};
############ END DEBUG ############*/
test_input[31464:31471] = '{32'hc19f697a, 32'hc1c071a1, 32'hc1641b70, 32'h4288c855, 32'hc2a3ebc1, 32'h42040ae1, 32'h427b7f7a, 32'hc22546fa};
test_label[3933] = '{32'hc22546fa};
test_output[3933] = '{32'h42db6ddf};
/*############ DEBUG ############
test_input[31464:31471] = '{-19.9265015988, -24.0554830812, -14.2566989596, 68.3912703064, -81.9604591524, 33.0106240247, 62.8744904664, -41.3193112343};
test_label[3933] = '{-41.3193112343};
test_output[3933] = '{109.714592255};
############ END DEBUG ############*/
test_input[31472:31479] = '{32'hc21b0018, 32'hbf9c1528, 32'hc267e64a, 32'h42265ed8, 32'hc288be40, 32'h4187d5dd, 32'h42a1fbe9, 32'h41dded58};
test_label[3934] = '{32'hc21b0018};
test_output[3934] = '{32'h42ef7bf5};
/*############ DEBUG ############
test_input[31472:31479] = '{-38.7500926269, -1.21939559683, -57.9748899179, 41.5926206627, -68.3715856375, 16.9794247346, 80.9920092636, 27.7408895871};
test_label[3934] = '{-38.7500926269};
test_output[3934] = '{119.742101891};
############ END DEBUG ############*/
test_input[31480:31487] = '{32'h40943ad7, 32'h414e54f5, 32'h42583be1, 32'hc289195d, 32'h423ae011, 32'hc2a29ec4, 32'hc2a23751, 32'h42810e48};
test_label[3935] = '{32'h40943ad7};
test_output[3935] = '{32'h426f953c};
/*############ DEBUG ############
test_input[31480:31487] = '{4.63218236954, 12.8957417771, 54.0584749954, -68.5495387824, 46.7188157039, -81.3100855588, -81.1080397168, 64.5278920352};
test_label[3935] = '{4.63218236954};
test_output[3935] = '{59.8957380753};
############ END DEBUG ############*/
test_input[31488:31495] = '{32'hc29b3916, 32'hc085b1b4, 32'hc29d25ce, 32'h4281fdf1, 32'h41d33b4c, 32'hc2c7ad5e, 32'hc276cc69, 32'hc1070c2c};
test_label[3936] = '{32'hc29d25ce};
test_output[3936] = '{32'h430f91e0};
/*############ DEBUG ############
test_input[31488:31495] = '{-77.6114958963, -4.17794240939, -78.5738407725, 64.9959811711, 26.4039543174, -99.8386054011, -61.6996184911, -8.44047192365};
test_label[3936] = '{-78.5738407725};
test_output[3936] = '{143.569821944};
############ END DEBUG ############*/
test_input[31496:31503] = '{32'h42823514, 32'hc2c1bf97, 32'hc254500c, 32'hc24fe429, 32'h429d55b5, 32'h40e5cffc, 32'hc125c7ff, 32'h42b301d2};
test_label[3937] = '{32'hc2c1bf97};
test_output[3937] = '{32'h433a60b6};
/*############ DEBUG ############
test_input[31496:31503] = '{65.1036715747, -96.8741994876, -53.0781722834, -51.9728140497, 78.6673958548, 7.18163853158, -10.3613271068, 89.5035581939};
test_label[3937] = '{-96.8741994876};
test_output[3937] = '{186.377777356};
############ END DEBUG ############*/
test_input[31504:31511] = '{32'h40c6b4a0, 32'hc0c6b52f, 32'hc12961d3, 32'h424fa253, 32'h4183b5a7, 32'hc0af8f4e, 32'hc2c17ac7, 32'hc288356e};
test_label[3938] = '{32'hc0c6b52f};
test_output[3938] = '{32'h426878f9};
/*############ DEBUG ############
test_input[31504:31511] = '{6.20954913869, -6.20961722998, -10.5863824761, 51.9085204351, 16.4636971373, -5.48624340976, -96.7398004162, -68.1043554222};
test_label[3938] = '{-6.20961722998};
test_output[3938] = '{58.1181376651};
############ END DEBUG ############*/
test_input[31512:31519] = '{32'h4220288b, 32'hc29dde7e, 32'h4224e49f, 32'hc29440dc, 32'hc2679b01, 32'h42c50ef4, 32'h41f9daaa, 32'h41c43764};
test_label[3939] = '{32'h41c43764};
test_output[3939] = '{32'h4294011b};
/*############ DEBUG ############
test_input[31512:31519] = '{40.039591588, -78.9345565538, 41.2232619585, -74.1266810045, -57.9013728234, 98.5292034501, 31.2317699351, 24.5270469025};
test_label[3939] = '{24.5270469025};
test_output[3939] = '{74.0021565476};
############ END DEBUG ############*/
test_input[31520:31527] = '{32'hc289cd90, 32'hc1aff430, 32'h42b2eb0e, 32'h3fa80fc1, 32'hc2178ad7, 32'h4282f5ac, 32'h42169408, 32'hc28d26d8};
test_label[3940] = '{32'hc1aff430};
test_output[3940] = '{32'h42dee81a};
/*############ DEBUG ############
test_input[31520:31527] = '{-68.9014872843, -21.9942322212, 89.4590913923, 1.31298081048, -37.8855869922, 65.4798268059, 37.6445621568, -70.5758629588};
test_label[3940] = '{-21.9942322212};
test_output[3940] = '{111.453323614};
############ END DEBUG ############*/
test_input[31528:31535] = '{32'hc28bfc4d, 32'h429f08fa, 32'hc221e941, 32'h42bafb10, 32'h4293b4a2, 32'hc2810752, 32'hc1b68c88, 32'h4230544d};
test_label[3941] = '{32'h4293b4a2};
test_output[3941] = '{32'h419d19b6};
/*############ DEBUG ############
test_input[31528:31535] = '{-69.9927747941, 79.517535161, -40.4777855763, 93.4903545939, 73.8528008531, -64.5142981213, -22.8186188983, 44.0823259047};
test_label[3941] = '{73.8528008531};
test_output[3941] = '{19.6375545982};
############ END DEBUG ############*/
test_input[31536:31543] = '{32'hc2671870, 32'h41c4b991, 32'hc2b832b6, 32'hc2a6ca23, 32'h42a83f72, 32'h429bcc32, 32'hc28da40a, 32'hc1831e55};
test_label[3942] = '{32'hc2671870};
test_output[3942] = '{32'h430de657};
/*############ DEBUG ############
test_input[31536:31543] = '{-57.7738647316, 24.5906095474, -92.0990458547, -83.3947983279, 84.1239160118, 77.8988166527, -70.8203857272, -16.3898114093};
test_label[3942] = '{-57.7738647316};
test_output[3942] = '{141.899757915};
############ END DEBUG ############*/
test_input[31544:31551] = '{32'h42c2ec0b, 32'h4223bd6f, 32'hc1b0f108, 32'h428b2444, 32'h427eea01, 32'h4223b268, 32'h40d8b337, 32'h426d7729};
test_label[3943] = '{32'h427eea01};
test_output[3943] = '{32'h4206ee14};
/*############ DEBUG ############
test_input[31544:31551] = '{97.4610198346, 40.9349940915, -22.1176910029, 69.5708323953, 63.7285207283, 40.9242243105, 6.77187664215, 59.3663674896};
test_label[3943] = '{63.7285207283};
test_output[3943] = '{33.7324991063};
############ END DEBUG ############*/
test_input[31552:31559] = '{32'h42bf458d, 32'hc2ba2b50, 32'hc2859895, 32'h4108b3e2, 32'h428ec27a, 32'h4239b3d5, 32'h4131c39d, 32'h42983d28};
test_label[3944] = '{32'h4108b3e2};
test_output[3944] = '{32'h42ae2f10};
/*############ DEBUG ############
test_input[31552:31559] = '{95.6358390874, -93.0845963615, -66.7980088446, 8.5439169294, 71.3798352499, 46.4256168499, 11.1102567855, 76.1194474402};
test_label[3944] = '{8.5439169294};
test_output[3944] = '{87.0919221613};
############ END DEBUG ############*/
test_input[31560:31567] = '{32'hc1e266a9, 32'h422863e6, 32'hc231a59b, 32'hc1233f2e, 32'hc20f6c22, 32'hc29bc6e2, 32'hc27670c4, 32'hc209809c};
test_label[3945] = '{32'hc27670c4};
test_output[3945] = '{32'h42cf6a55};
/*############ DEBUG ############
test_input[31560:31567] = '{-28.3001274566, 42.0975573555, -44.4117247379, -10.2029248735, -35.8555980854, -77.8884396776, -61.6101226769, -34.3755933967};
test_label[3945] = '{-61.6101226769};
test_output[3945] = '{103.707680032};
############ END DEBUG ############*/
test_input[31568:31575] = '{32'hc1e274ad, 32'h42a34998, 32'h421d4c55, 32'hc12cd5ba, 32'hc2ab6f8d, 32'hc1f22384, 32'h4287a8b1, 32'hc28c75b8};
test_label[3946] = '{32'hc1f22384};
test_output[3946] = '{32'h42dfd279};
/*############ DEBUG ############
test_input[31568:31575] = '{-28.3069700279, 81.6437347661, 39.3245439429, -10.8021791781, -85.7178705767, -30.2673416055, 67.8294791811, -70.2299200954};
test_label[3946] = '{-30.2673416055};
test_output[3946] = '{111.911077373};
############ END DEBUG ############*/
test_input[31576:31583] = '{32'h41d698e0, 32'h42c159c3, 32'h42c79028, 32'hc2b9f064, 32'h3f8a1a0d, 32'h42b755bc, 32'hc2688dce, 32'h428228e8};
test_label[3947] = '{32'h3f8a1a0d};
test_output[3947] = '{32'h42c57e52};
/*############ DEBUG ############
test_input[31576:31583] = '{26.8246464093, 96.6753171044, 99.781555471, -92.9695149496, 1.07891998948, 91.667447442, -58.1384797039, 65.0798984465};
test_label[3947] = '{1.07891998948};
test_output[3947] = '{98.746717753};
############ END DEBUG ############*/
test_input[31584:31591] = '{32'hc0281a1c, 32'h429959fb, 32'hc2a90d15, 32'hc22de8d5, 32'hc2974969, 32'hc1589b66, 32'hc2c094fd, 32'h41f393f6};
test_label[3948] = '{32'hc2a90d15};
test_output[3948] = '{32'h43213388};
/*############ DEBUG ############
test_input[31584:31591] = '{-2.62659357554, 76.6757407106, -84.5255532292, -43.4773751719, -75.6433781299, -13.5379395405, -96.2909902878, 30.4472464046};
test_label[3948] = '{-84.5255532292};
test_output[3948] = '{161.20129394};
############ END DEBUG ############*/
test_input[31592:31599] = '{32'hc1dc980d, 32'h417ae96c, 32'hc22b540c, 32'h40171165, 32'hc241d6f2, 32'h41ddf8ef, 32'hc291872c, 32'hc2b7ee21};
test_label[3949] = '{32'hc291872c};
test_output[3949] = '{32'h42c90569};
/*############ DEBUG ############
test_input[31592:31599] = '{-27.5742428098, 15.6819874476, -42.8320781362, 2.36043675369, -48.459907587, 27.7465500957, -72.7640098814, -91.9650919129};
test_label[3949] = '{-72.7640098814};
test_output[3949] = '{100.510565737};
############ END DEBUG ############*/
test_input[31600:31607] = '{32'h42bc4619, 32'h41bf9ecc, 32'hc21686a5, 32'h41f62c6c, 32'h42163033, 32'hc2bd7a28, 32'hc24dfd0e, 32'h42b5a2a3};
test_label[3950] = '{32'hc21686a5};
test_output[3950] = '{32'h4303cdcf};
/*############ DEBUG ############
test_input[31600:31607] = '{94.1369098791, 23.9525374531, -37.6314900103, 30.7716907762, 37.5470689912, -94.7385862592, -51.4971237744, 90.8176522047};
test_label[3950] = '{-37.6314900103};
test_output[3950] = '{131.803940453};
############ END DEBUG ############*/
test_input[31608:31615] = '{32'h41fb0d0d, 32'hc2a36c5f, 32'hc29b8f49, 32'hc18058e9, 32'h428b3195, 32'hc205a6bf, 32'h3fb9782e, 32'hc13ef852};
test_label[3951] = '{32'hc18058e9};
test_output[3951] = '{32'h42ab47cf};
/*############ DEBUG ############
test_input[31608:31615] = '{31.3813719138, -81.711659137, -77.7798516177, -16.0434140812, 69.5968403608, -33.4128395435, 1.44898003409, -11.9356253164};
test_label[3951] = '{-16.0434140812};
test_output[3951] = '{85.640254442};
############ END DEBUG ############*/
test_input[31616:31623] = '{32'h42ba4974, 32'h42600a33, 32'hc28e8813, 32'hc2c2817d, 32'hc233d542, 32'hc1ed4254, 32'h424c626a, 32'h42ab811a};
test_label[3952] = '{32'h42ba4974};
test_output[3952] = '{32'h3a2195ac};
/*############ DEBUG ############
test_input[31616:31623] = '{93.1434633665, 56.0099609493, -71.2657710176, -97.25290956, -44.9582593999, -29.6573872458, 51.0961059204, 85.752151557};
test_label[3952] = '{93.1434633665};
test_output[3952] = '{0.000616396567258};
############ END DEBUG ############*/
test_input[31624:31631] = '{32'hc29275be, 32'hc13dc037, 32'h4289dfb9, 32'hc2abfdbf, 32'h41ffb412, 32'h42b8e12a, 32'h42b258f7, 32'hc20e7243};
test_label[3953] = '{32'h4289dfb9};
test_output[3953] = '{32'h41bc5275};
/*############ DEBUG ############
test_input[31624:31631] = '{-73.2299676065, -11.8594271321, 68.9369592622, -85.9956001726, 31.9629244713, 92.4397734319, 89.1737599181, -35.61158344};
test_label[3953] = '{68.9369592622};
test_output[3953] = '{23.5402623914};
############ END DEBUG ############*/
test_input[31632:31639] = '{32'h4245c984, 32'h428addb7, 32'h42a7c91a, 32'hc27cd95c, 32'hc25c2702, 32'hc29f2e06, 32'hc1f0b5db, 32'h40ff2887};
test_label[3954] = '{32'hc29f2e06};
test_output[3954] = '{32'h43237b90};
/*############ DEBUG ############
test_input[31632:31639] = '{49.4467920611, 69.4330377452, 83.892775263, -63.2122631714, -55.0380934118, -79.5898878806, -30.0887962481, 7.97369708405};
test_label[3954] = '{-79.5898878806};
test_output[3954] = '{163.482663669};
############ END DEBUG ############*/
test_input[31640:31647] = '{32'hc23c12a8, 32'h4284e37e, 32'h416e36db, 32'hc2208019, 32'hc2996ff7, 32'hbf6947e0, 32'h429680bd, 32'hc1bac32e};
test_label[3955] = '{32'hc2208019};
test_output[3955] = '{32'h42e6c0dd};
/*############ DEBUG ############
test_input[31640:31647] = '{-47.0182178026, 66.4443173393, 14.8883921841, -40.125096361, -76.7186782436, -0.911253003646, 75.2514427519, -23.345303459};
test_label[3955] = '{-40.125096361};
test_output[3955] = '{115.376688765};
############ END DEBUG ############*/
test_input[31648:31655] = '{32'hc2a86e95, 32'hc28c3210, 32'h422b3bf8, 32'h42b7b874, 32'hc2ab114b, 32'hc2b1a30b, 32'hc285171d, 32'h405713d1};
test_label[3956] = '{32'hc28c3210};
test_output[3956] = '{32'h4321f542};
/*############ DEBUG ############
test_input[31648:31655] = '{-84.2159774806, -70.0977764978, 42.8085622853, 91.8602580248, -85.5337730902, -88.8184465392, -66.5451449254, 3.36058459324};
test_label[3956] = '{-70.0977764978};
test_output[3956] = '{161.958034523};
############ END DEBUG ############*/
test_input[31656:31663] = '{32'hc1a590b3, 32'h4260f0ec, 32'h41732c1d, 32'h42c24a83, 32'hc272126d, 32'hc22d8ca9, 32'hc0b7b26a, 32'h42783b23};
test_label[3957] = '{32'hc22d8ca9};
test_output[3957] = '{32'h430c886c};
/*############ DEBUG ############
test_input[31656:31663] = '{-20.6956530917, 56.2352753142, 15.1982694964, 97.1455289901, -60.5179949693, -43.3873635689, -5.74052902317, 62.057749312};
test_label[3957] = '{-43.3873635689};
test_output[3957] = '{140.532892559};
############ END DEBUG ############*/
test_input[31664:31671] = '{32'hc1a253cc, 32'hc2954c41, 32'hc1a040e2, 32'h41f135cd, 32'h40068b5c, 32'h42a30f7d, 32'h4242850f, 32'hc1ae0b59};
test_label[3958] = '{32'hc2954c41};
test_output[3958] = '{32'h431c2ddf};
/*############ DEBUG ############
test_input[31664:31671] = '{-20.2909169991, -74.6489352343, -20.0316805587, 30.1512702309, 2.10225573632, 81.530252449, 48.629940849, -21.7555415792};
test_label[3958] = '{-74.6489352343};
test_output[3958] = '{156.179187683};
############ END DEBUG ############*/
test_input[31672:31679] = '{32'h4294459e, 32'hc22ea618, 32'hc19aaaeb, 32'h4295b3a9, 32'hc13182d8, 32'hc2bc1bb4, 32'hbf8c83a3, 32'h4231b19e};
test_label[3959] = '{32'hc2bc1bb4};
test_output[3959] = '{32'h43294da3};
/*############ DEBUG ############
test_input[31672:31679] = '{74.1359733444, -43.6622017085, -19.3334551246, 74.8509008525, -11.0944443963, -94.0541078527, -1.09776726057, 44.4234531299};
test_label[3959] = '{-94.0541078527};
test_output[3959] = '{169.303266285};
############ END DEBUG ############*/
test_input[31680:31687] = '{32'hc24bb23c, 32'h4237ca7e, 32'h41ab25bc, 32'hc1f5c3c3, 32'hc1b9498f, 32'h42a7818c, 32'hc2bde1e7, 32'hc2820a16};
test_label[3960] = '{32'hc2820a16};
test_output[3960] = '{32'h4314c5d1};
/*############ DEBUG ############
test_input[31680:31687] = '{-50.9240551735, 45.9477461644, 21.3934246689, -30.7205862767, -23.1609176805, 83.7530240638, -94.9412182175, -65.0197014766};
test_label[3960] = '{-65.0197014766};
test_output[3960] = '{148.77272554};
############ END DEBUG ############*/
test_input[31688:31695] = '{32'h42995da6, 32'h418f4db3, 32'h4206df47, 32'h42c6b8c4, 32'hc1549e43, 32'hc2acda64, 32'hc235094b, 32'h42c44498};
test_label[3961] = '{32'h42995da6};
test_output[3961] = '{32'h41b77b10};
/*############ DEBUG ############
test_input[31688:31695] = '{76.6829048355, 17.9129395878, 33.7180451477, 99.3608738667, -13.2886384608, -86.4265430788, -45.2590744844, 98.1339728845};
test_label[3961] = '{76.6829048355};
test_output[3961] = '{22.9350886455};
############ END DEBUG ############*/
test_input[31696:31703] = '{32'h42b40587, 32'h421881d6, 32'hc2656a9e, 32'hc2af5f04, 32'h4236207d, 32'hc136d672, 32'h42a9c8a4, 32'hc22e0455};
test_label[3962] = '{32'h4236207d};
test_output[3962] = '{32'h4231f0ac};
/*############ DEBUG ############
test_input[31696:31703] = '{90.01079468, 38.1267945596, -57.3541193614, -87.6855789525, 45.5317283522, -11.4273550852, 84.8918766304, -43.5042308876};
test_label[3962] = '{45.5317283522};
test_output[3962] = '{44.4850309959};
############ END DEBUG ############*/
test_input[31704:31711] = '{32'hc264b143, 32'h42b59d4f, 32'hc2608621, 32'hc1067d23, 32'h42a6e5f2, 32'h419baeb0, 32'h42351fbe, 32'h428b8fbd};
test_label[3963] = '{32'h42b59d4f};
test_output[3963] = '{32'h3a2708c8};
/*############ DEBUG ############
test_input[31704:31711] = '{-57.173106308, 90.8072412669, -56.1309852983, -8.40555106793, 83.4491086872, 19.4602971557, 45.2809971225, 69.7807388693};
test_label[3963] = '{90.8072412669};
test_output[3963] = '{0.000637185312164};
############ END DEBUG ############*/
test_input[31712:31719] = '{32'h41aae469, 32'h42bc4c2f, 32'h40ecb5ed, 32'h40a8fdea, 32'hc18ae7a8, 32'hc1c8bf39, 32'hc0af62cf, 32'hc0a1ce8f};
test_label[3964] = '{32'hc0a1ce8f};
test_output[3964] = '{32'h42c66918};
/*############ DEBUG ############
test_input[31712:31719] = '{21.3615283764, 94.1487939264, 7.39720795944, 5.28099528294, -17.363113454, -25.0933708913, -5.48081151431, -5.05646453101};
test_label[3964] = '{-5.05646453101};
test_output[3964] = '{99.2052584574};
############ END DEBUG ############*/
test_input[31720:31727] = '{32'hc204bfb4, 32'h428173b8, 32'hc2aec3fd, 32'h415a09fe, 32'h416b7b21, 32'hc2b8b9be, 32'h41c89a07, 32'hc24bd8ec};
test_label[3965] = '{32'hc2aec3fd};
test_output[3965] = '{32'h43181bdb};
/*############ DEBUG ############
test_input[31720:31727] = '{-33.1872115796, 64.7260120872, -87.3827918561, 13.6274395945, 14.7175611052, -92.3627804253, 25.0752087074, -50.9618369371};
test_label[3965] = '{-87.3827918561};
test_output[3965] = '{152.108803943};
############ END DEBUG ############*/
test_input[31728:31735] = '{32'h42871f0a, 32'hc1f2297e, 32'h42c5a8ec, 32'h427eb4d7, 32'h40912260, 32'h4243c0fd, 32'hc2b40230, 32'hc27df933};
test_label[3966] = '{32'h42c5a8ec};
test_output[3966] = '{32'h28f20000};
/*############ DEBUG ############
test_input[31728:31735] = '{67.5606224226, -30.2702596905, 98.8299291465, 63.6766032019, 4.53544632503, 48.938464191, -90.0042734246, -63.4933579858};
test_label[3966] = '{98.8299291465};
test_output[3966] = '{2.68673971959e-14};
############ END DEBUG ############*/
test_input[31736:31743] = '{32'hc2b04d0a, 32'hc243f603, 32'hc0fa9774, 32'h412013dc, 32'hc1cda490, 32'h4287ec0d, 32'hc2b410e9, 32'hc1f64c9d};
test_label[3967] = '{32'hc2b04d0a};
test_output[3967] = '{32'h431c1c8c};
/*############ DEBUG ############
test_input[31736:31743] = '{-88.1504691731, -48.9902472667, -7.83098798558, 10.0048488913, -25.7053535864, 67.9610389695, -90.0330278445, -30.7874097347};
test_label[3967] = '{-88.1504691731};
test_output[3967] = '{156.111508143};
############ END DEBUG ############*/
test_input[31744:31751] = '{32'hc2b05d29, 32'hc260f0d5, 32'hc240ae4a, 32'h4074083e, 32'h4212839f, 32'hc12e5eb7, 32'hc2ae0a35, 32'h42bcea70};
test_label[3968] = '{32'hc2ae0a35};
test_output[3968] = '{32'h43357a53};
/*############ DEBUG ############
test_input[31744:31751] = '{-88.1819569795, -56.2351883587, -48.1702050688, 3.81300311258, 36.6285374579, -10.8981238647, -87.0199370176, 94.4578868745};
test_label[3968] = '{-87.0199370176};
test_output[3968] = '{181.477823892};
############ END DEBUG ############*/
test_input[31752:31759] = '{32'hc14119a2, 32'h42ae0747, 32'h42c30303, 32'h4296c074, 32'h42a5fdc1, 32'h4255bd2f, 32'h4215daf7, 32'h4287c6ad};
test_label[3969] = '{32'h4215daf7};
test_output[3969] = '{32'h42702b16};
/*############ DEBUG ############
test_input[31752:31759] = '{-12.0687580871, 87.0142124563, 97.5058797418, 75.3758882619, 82.9956146365, 53.4347494428, 37.4638333631, 67.8880382786};
test_label[3969] = '{37.4638333631};
test_output[3969] = '{60.0420746446};
############ END DEBUG ############*/
test_input[31760:31767] = '{32'hc21fe621, 32'h424ad0e1, 32'h41c5c100, 32'hc13020ea, 32'h424a448d, 32'h42acebdb, 32'h42b84b65, 32'hc262ae01};
test_label[3970] = '{32'h41c5c100};
test_output[3970] = '{32'h4286dce1};
/*############ DEBUG ############
test_input[31760:31767] = '{-39.9747343822, 50.7039847971, 24.7192378946, -11.0080355062, 50.5669455139, 86.4606555134, 92.1472573297, -56.6699259474};
test_label[3970] = '{24.7192378946};
test_output[3970] = '{67.4314047952};
############ END DEBUG ############*/
test_input[31768:31775] = '{32'h4271b1c7, 32'hc2301217, 32'h42472f59, 32'hc2c4edcf, 32'hc2984d4f, 32'hbfd76fb3, 32'h41612c2a, 32'hc2af312e};
test_label[3971] = '{32'h41612c2a};
test_output[3971] = '{32'h423966c3};
/*############ DEBUG ############
test_input[31768:31775] = '{60.4236102838, -44.0176662418, 49.7962361569, -98.46447063, -76.1509948605, -1.68309632421, 14.0732821122, -87.5960556477};
test_label[3971] = '{14.0732821122};
test_output[3971] = '{46.3503524146};
############ END DEBUG ############*/
test_input[31776:31783] = '{32'hc2b6509e, 32'hc2968ee1, 32'hc2183e56, 32'h41bd849b, 32'h429eb7bb, 32'hc2604f9c, 32'h420497f8, 32'h428b2842};
test_label[3972] = '{32'hc2968ee1};
test_output[3972] = '{32'h431aa352};
/*############ DEBUG ############
test_input[31776:31783] = '{-91.1574516964, -75.2790603843, -38.0608740813, 23.6897484888, 79.3588521073, -56.0777420513, 33.148408068, 69.5786277575};
test_label[3972] = '{-75.2790603843};
test_output[3972] = '{154.637969049};
############ END DEBUG ############*/
test_input[31784:31791] = '{32'h42784219, 32'hc28bd0e2, 32'h40881c37, 32'h4290866a, 32'hc2a1730f, 32'hc2c20fa4, 32'hc2baaa4a, 32'h429b3877};
test_label[3973] = '{32'hc28bd0e2};
test_output[3973] = '{32'h431385e4};
/*############ DEBUG ############
test_input[31784:31791] = '{62.064548918, -69.9079772263, 4.25344442512, 72.2625299058, -80.724723888, -97.030550057, -93.3325937483, 77.6102804854};
test_label[3973] = '{-69.9079772263};
test_output[3973] = '{147.523005444};
############ END DEBUG ############*/
test_input[31792:31799] = '{32'h418cd33d, 32'hc25c7541, 32'hc2844b61, 32'hc2c153e2, 32'h41d1ee61, 32'hc2b6b63a, 32'h42c3ee95, 32'h41718b62};
test_label[3974] = '{32'h42c3ee95};
test_output[3974] = '{32'h80000000};
/*############ DEBUG ############
test_input[31792:31799] = '{17.6031445539, -55.1145065643, -66.1472245069, -96.6638329732, 26.24139634, -91.3559087226, 97.9659802644, 15.0965292545};
test_label[3974] = '{97.9659802644};
test_output[3974] = '{-0.0};
############ END DEBUG ############*/
test_input[31800:31807] = '{32'hbf345d96, 32'hc297e086, 32'hc22dea60, 32'hc27bd2d4, 32'hc293cfd4, 32'hc2b1b836, 32'hc210d148, 32'h42bdde59};
test_label[3975] = '{32'hc210d148};
test_output[3975] = '{32'h4303237f};
/*############ DEBUG ############
test_input[31800:31807] = '{-0.704553036034, -75.9385195634, -43.4788809085, -62.9558881641, -73.9059131981, -88.8597893307, -36.2043767905, 94.9342723251};
test_label[3975] = '{-36.2043767905};
test_output[3975] = '{131.138649116};
############ END DEBUG ############*/
test_input[31808:31815] = '{32'h42a4b308, 32'h4280b4fd, 32'h4216d67d, 32'h4296a8f0, 32'h419e912b, 32'h429ceb5a, 32'hc1036d66, 32'hc26ef1df};
test_label[3976] = '{32'h4280b4fd};
test_output[3976] = '{32'h41902369};
/*############ DEBUG ############
test_input[31808:31815] = '{82.3496672735, 64.3534921604, 37.7094630545, 75.3299545083, 19.8208820243, 78.459669727, -8.21420820319, -59.7362018051};
test_label[3976] = '{64.3534921604};
test_output[3976] = '{18.0172901081};
############ END DEBUG ############*/
test_input[31816:31823] = '{32'h4109b9f6, 32'h42c60771, 32'hc21270f0, 32'h4260d126, 32'hc24a3a5a, 32'hc22b7279, 32'h421f7f5b, 32'h41fa30cc};
test_label[3977] = '{32'h42c60771};
test_output[3977] = '{32'h80000000};
/*############ DEBUG ############
test_input[31816:31823] = '{8.60790051693, 99.0145306485, -36.6102903514, 56.2042472578, -50.5569839773, -42.8617878362, 39.8743713891, 31.2738267287};
test_label[3977] = '{99.0145306485};
test_output[3977] = '{-0.0};
############ END DEBUG ############*/
test_input[31824:31831] = '{32'h419ab75f, 32'hc2b71708, 32'hc1d4d7a6, 32'hc2472ad6, 32'hc2523312, 32'hc2a67e15, 32'hc130d519, 32'hc27be7b2};
test_label[3978] = '{32'hc2a67e15};
test_output[3978] = '{32'h42cd2bed};
/*############ DEBUG ############
test_input[31824:31831] = '{19.3395362179, -91.544981258, -26.6052968541, -49.7918331106, -52.5498750874, -83.2462533412, -11.052026006, -62.9762655301};
test_label[3978] = '{-83.2462533412};
test_output[3978] = '{102.585789559};
############ END DEBUG ############*/
test_input[31832:31839] = '{32'h429f784b, 32'hc2109bd5, 32'hc1efd5f7, 32'h427cef9b, 32'h4119adf9, 32'hc22dfca2, 32'h4262eda5, 32'hc203cb9a};
test_label[3979] = '{32'hc203cb9a};
test_output[3979] = '{32'h42e15e18};
/*############ DEBUG ############
test_input[31832:31839] = '{79.7349462841, -36.1521784175, -29.9794747033, 63.2339882695, 9.604973999, -43.4967098696, 56.7320750341, -32.9488300031};
test_label[3979] = '{-32.9488300031};
test_output[3979] = '{112.683776355};
############ END DEBUG ############*/
test_input[31840:31847] = '{32'h41a913c0, 32'h41cb084e, 32'hc2552ecf, 32'h3f414a3e, 32'h42ac96d0, 32'h429072cd, 32'h4267cfee, 32'hc2918440};
test_label[3980] = '{32'h4267cfee};
test_output[3980] = '{32'h41e2bb64};
/*############ DEBUG ############
test_input[31840:31847] = '{21.1346427439, 25.3790546938, -53.2957127272, 0.755039104012, 86.2945544072, 72.2242188454, 57.9530562987, -72.7582994585};
test_label[3980] = '{57.9530562987};
test_output[3980] = '{28.3414988835};
############ END DEBUG ############*/
test_input[31848:31855] = '{32'hc2369970, 32'hbef771fe, 32'h41a2ca9b, 32'h42b4e276, 32'hc0cd3ce7, 32'hc22eee22, 32'hc26e6ee3, 32'hc201dbc7};
test_label[3981] = '{32'h42b4e276};
test_output[3981] = '{32'h80000000};
/*############ DEBUG ############
test_input[31848:31855] = '{-45.6498403616, -0.483291566963, 20.3489290085, 90.4423070165, -6.41368436773, -43.7325513591, -59.6082868292, -32.464628128};
test_label[3981] = '{90.4423070165};
test_output[3981] = '{-0.0};
############ END DEBUG ############*/
test_input[31856:31863] = '{32'h42bf25ec, 32'h42b60caa, 32'hc200a2a1, 32'hc2a9faf4, 32'h41d992d3, 32'hc236874e, 32'hc2405b02, 32'hc2234585};
test_label[3982] = '{32'hc200a2a1};
test_output[3982] = '{32'h42ff7ca0};
/*############ DEBUG ############
test_input[31856:31863] = '{95.5740698206, 91.024731375, -32.1588165345, -84.9901464132, 27.1966922267, -45.6321337695, -48.0888739879, -40.8178912256};
test_label[3982] = '{-32.1588165345};
test_output[3982] = '{127.743405037};
############ END DEBUG ############*/
test_input[31864:31871] = '{32'hc1ce1559, 32'h4193a4f0, 32'h4230bf0a, 32'h424fef3c, 32'h40c8fe7e, 32'hc1f6841e, 32'h41018731, 32'hc110179c};
test_label[3983] = '{32'hc1ce1559};
test_output[3983] = '{32'h429b7d2a};
/*############ DEBUG ############
test_input[31864:31871] = '{-25.7604244926, 18.4555358908, 44.1865628562, 51.9836273677, 6.28106609382, -30.814511034, 8.09550536365, -9.00576399649};
test_label[3983] = '{-25.7604244926};
test_output[3983] = '{77.7444627154};
############ END DEBUG ############*/
test_input[31872:31879] = '{32'h41b19a3a, 32'hc248ce6a, 32'hc1c80349, 32'hc283583a, 32'hc2c471d6, 32'h4232ddd1, 32'h42b55565, 32'hc1ce75af};
test_label[3984] = '{32'hc2c471d6};
test_output[3984] = '{32'h433ce39d};
/*############ DEBUG ############
test_input[31872:31879] = '{22.2003051481, -50.2015764404, -25.0016043344, -65.6723205518, -98.2223323946, 44.7166178319, 90.6667883259, -25.8074621937};
test_label[3984] = '{-98.2223323946};
test_output[3984] = '{188.88912072};
############ END DEBUG ############*/
test_input[31880:31887] = '{32'h429c8858, 32'hc21f3038, 32'h427cfb00, 32'h42b9a0ff, 32'hc2471e20, 32'hc23ae9c0, 32'hc2a6e706, 32'hc295e331};
test_label[3985] = '{32'hc23ae9c0};
test_output[3985] = '{32'h430b8aef};
/*############ DEBUG ############
test_input[31880:31887] = '{78.2662952663, -39.7970874893, 63.245116799, 92.8144423607, -49.779417182, -46.7282700469, -83.451219646, -74.9437313883};
test_label[3985] = '{-46.7282700469};
test_output[3985] = '{139.542712888};
############ END DEBUG ############*/
test_input[31888:31895] = '{32'h420f698f, 32'h41832d0d, 32'hc29572a7, 32'h41b73474, 32'h41ccce83, 32'hc01e4654, 32'h428ee232, 32'hc110770c};
test_label[3986] = '{32'h41b73474};
test_output[3986] = '{32'h42422a2b};
/*############ DEBUG ############
test_input[31888:31895] = '{35.8530832075, 16.3969982111, -74.7239289624, 22.9006122382, 25.6008355531, -2.4730425278, 71.4417912332, -9.02906397117};
test_label[3986] = '{22.9006122382};
test_output[3986] = '{48.541178995};
############ END DEBUG ############*/
test_input[31896:31903] = '{32'hc2ace5b9, 32'h41e995e7, 32'hc2b90c08, 32'h41f3a59b, 32'h4254de24, 32'h419f1d4b, 32'hc204f023, 32'h42ae01ea};
test_label[3987] = '{32'h41f3a59b};
test_output[3987] = '{32'h42623106};
/*############ DEBUG ############
test_input[31896:31903] = '{-86.4486765452, 29.198195182, -92.5235017, 30.4558615171, 53.2169360331, 19.8893040277, -33.2345098241, 87.0037353028};
test_label[3987] = '{30.4558615171};
test_output[3987] = '{56.5478737857};
############ END DEBUG ############*/
test_input[31904:31911] = '{32'h411d898b, 32'hc23c2efa, 32'hc29c78a2, 32'hc20264fe, 32'hc1bf0c74, 32'h41b13a39, 32'hc244f867, 32'hc22abc2a};
test_label[3988] = '{32'hc244f867};
test_output[3988] = '{32'h428ecac2};
/*############ DEBUG ############
test_input[31904:31911] = '{9.84607953079, -47.0458742419, -78.2356118007, -32.5986262086, -23.881081211, 22.1534290468, -49.2425815815, -42.6837538735};
test_label[3988] = '{-49.2425815815};
test_output[3988] = '{71.3960151467};
############ END DEBUG ############*/
test_input[31912:31919] = '{32'h414bec39, 32'h42495669, 32'h429d62d5, 32'hc286a18a, 32'hc256d573, 32'hc13d7712, 32'h41a0da9d, 32'hc252d051};
test_label[3989] = '{32'hc13d7712};
test_output[3989] = '{32'h42b511b7};
/*############ DEBUG ############
test_input[31912:31919] = '{12.74517111, 50.3343852934, 78.6930293848, -67.3155097593, -53.708446849, -11.8415698947, 20.1067450207, -52.7034344288};
test_label[3989] = '{-11.8415698947};
test_output[3989] = '{90.5345992795};
############ END DEBUG ############*/
test_input[31920:31927] = '{32'hc242364c, 32'h41129bc0, 32'hc2695078, 32'hc27ada21, 32'h42bd663a, 32'h42b9e230, 32'hc2a5cd90, 32'hc1c714d7};
test_label[3990] = '{32'h42b9e230};
test_output[3990] = '{32'h3ff55e90};
/*############ DEBUG ############
test_input[31920:31927] = '{-48.5530244651, 9.1630248767, -58.3285843602, -62.7130157229, 94.6996643413, 92.9417762389, -82.9014884921, -24.885174912};
test_label[3990] = '{92.9417762389};
test_output[3990] = '{1.91694835808};
############ END DEBUG ############*/
test_input[31928:31935] = '{32'hc1c91c98, 32'h42566845, 32'hc162b966, 32'h426c6f0d, 32'hc2c6b1a3, 32'h4288845f, 32'hc109c3dd, 32'h417ed478};
test_label[3991] = '{32'h42566845};
test_output[3991] = '{32'h416a8251};
/*############ DEBUG ############
test_input[31928:31935] = '{-25.1389618, 53.6018264042, -14.1702633506, 59.108446857, -99.3469479344, 68.2585350173, -8.6103184802, 15.9268721968};
test_label[3991] = '{53.6018264042};
test_output[3991] = '{14.656815249};
############ END DEBUG ############*/
test_input[31936:31943] = '{32'hc031b020, 32'h42905015, 32'h422cd22c, 32'h4001d557, 32'hc2bd5bda, 32'h42a583e1, 32'h40ffc84a, 32'h422bf4bb};
test_label[3992] = '{32'h422bf4bb};
test_output[3992] = '{32'h421f130d};
/*############ DEBUG ############
test_input[31936:31943] = '{-2.77637485759, 72.1564065857, 43.205246563, 2.02864631996, -94.6793980298, 82.7575758377, 7.99319951202, 42.9889953815};
test_label[3992] = '{42.9889953815};
test_output[3992] = '{39.7686053428};
############ END DEBUG ############*/
test_input[31944:31951] = '{32'h42b4edf5, 32'hc24d3faa, 32'h42887dd6, 32'h42c0d811, 32'hc29bcfa8, 32'h42b7bcd2, 32'h4285ae5a, 32'hc1fa9cd4};
test_label[3993] = '{32'h42b7bcd2};
test_output[3993] = '{32'h40921eb7};
/*############ DEBUG ############
test_input[31944:31951] = '{90.4647599013, -51.3121736419, 68.2457697661, 96.4220049068, -77.905576027, 91.8687906476, 66.8405294631, -31.3265759611};
test_label[3993] = '{91.8687906476};
test_output[3993] = '{4.56624925588};
############ END DEBUG ############*/
test_input[31952:31959] = '{32'hc10d93dd, 32'h4039b3eb, 32'h41d68f76, 32'h4201e0e2, 32'h41fded19, 32'hc2687645, 32'hc2911bc6, 32'hc292eaa3};
test_label[3994] = '{32'h4039b3eb};
test_output[3994] = '{32'h41efb672};
/*############ DEBUG ############
test_input[31952:31959] = '{-8.84859979971, 2.90160629016, 26.8200499713, 32.469613463, 31.7407697267, -58.1154986716, -72.5542466664, -73.4582781101};
test_label[3994] = '{2.90160629016};
test_output[3994] = '{29.9640854144};
############ END DEBUG ############*/
test_input[31960:31967] = '{32'hc197720f, 32'hc17ecfff, 32'h422b6fd4, 32'hc24f55e6, 32'hc2ba7e70, 32'h42ac3ca6, 32'hc25558ee, 32'hc1630921};
test_label[3995] = '{32'hc1630921};
test_output[3995] = '{32'h42c89dca};
/*############ DEBUG ############
test_input[31960:31967] = '{-18.9306930976, -15.9257801806, 42.859206952, -51.8338868275, -93.2469481673, 86.1184527242, -53.3368465574, -14.1897287388};
test_label[3995] = '{-14.1897287388};
test_output[3995] = '{100.308181463};
############ END DEBUG ############*/
test_input[31968:31975] = '{32'hc25ac6db, 32'hc2411e5f, 32'h423234a8, 32'h42881b16, 32'hc22eebc6, 32'h422ab66e, 32'h42410b93, 32'hc2ad1f22};
test_label[3996] = '{32'hc2ad1f22};
test_output[3996] = '{32'h431a9d1c};
/*############ DEBUG ############
test_input[31968:31975] = '{-54.6941963121, -48.279658648, 44.5514207317, 68.0528989804, -43.7302466537, 42.6781524278, 48.2613028639, -86.5608091791};
test_label[3996] = '{-86.5608091791};
test_output[3996] = '{154.613708162};
############ END DEBUG ############*/
test_input[31976:31983] = '{32'h4112c160, 32'hbfe8c65e, 32'h428b4fab, 32'h41a47c67, 32'hc21b218c, 32'hc2818ee7, 32'h428d24cc, 32'h42a5e1b3};
test_label[3997] = '{32'h4112c160};
test_output[3997] = '{32'h42938988};
/*############ DEBUG ############
test_input[31976:31983] = '{9.17221070997, -1.81855374359, 69.6556001301, 20.5607437991, -38.7827608757, -64.7791089605, 70.5718687485, 82.9408184659};
test_label[3997] = '{9.17221070997};
test_output[3997] = '{73.7686137038};
############ END DEBUG ############*/
test_input[31984:31991] = '{32'hc2ba4965, 32'h424f1dd6, 32'h4101d25c, 32'hbf944cd3, 32'h41ae59d3, 32'hc29ca0e9, 32'hc1a2af48, 32'hc1e48332};
test_label[3998] = '{32'h424f1dd6};
test_output[3998] = '{32'h29d5c000};
/*############ DEBUG ############
test_input[31984:31991] = '{-93.1433451363, 51.7791373158, 8.11385751645, -1.15859447296, 21.7938589382, -78.3142803068, -20.3355866247, -28.5640601313};
test_label[3998] = '{51.7791373158};
test_output[3998] = '{9.49240686055e-14};
############ END DEBUG ############*/
test_input[31992:31999] = '{32'hc2be262e, 32'hc2bd331a, 32'hc258a710, 32'hc23e7f4a, 32'h40ca5f28, 32'hc2b95506, 32'hc1972894, 32'hc216bfa0};
test_label[3999] = '{32'hc2be262e};
test_output[3999] = '{32'h42cacc20};
/*############ DEBUG ############
test_input[31992:31999] = '{-95.0745673288, -94.5998076695, -54.1631459738, -47.624307048, 6.32411595204, -92.6660647269, -18.8948127086, -37.6871326935};
test_label[3999] = '{-95.0745673288};
test_output[3999] = '{101.398683281};
############ END DEBUG ############*/
test_input[32000:32007] = '{32'h4111b35f, 32'hc20fbf9e, 32'hc24ce5e0, 32'h40b0a937, 32'h41cfbac1, 32'h41a25777, 32'h41c60b1c, 32'h42bee0b7};
test_label[4000] = '{32'h40b0a937};
test_output[4000] = '{32'h42b3d624};
/*############ DEBUG ############
test_input[32000:32007] = '{9.10629207674, -35.9371262446, -51.2244884413, 5.52065614256, 25.9661893027, 20.2927081903, 24.7554253662, 95.4388986012};
test_label[4000] = '{5.52065614256};
test_output[4000] = '{89.9182424587};
############ END DEBUG ############*/
test_input[32008:32015] = '{32'hc2699fee, 32'h42bdc864, 32'hc174d12a, 32'h41a57dc5, 32'h427c7a56, 32'hc2c1a77b, 32'h423afed2, 32'hc0fceab2};
test_label[4001] = '{32'hc174d12a};
test_output[4001] = '{32'h42dc6289};
/*############ DEBUG ############
test_input[32008:32015] = '{-58.4061808763, 94.8913881826, -15.3010654772, 20.6864106845, 63.1194700287, -96.8271069302, 46.7488466647, -7.90364949395};
test_label[4001] = '{-15.3010654772};
test_output[4001] = '{110.19245366};
############ END DEBUG ############*/
test_input[32016:32023] = '{32'h4296601c, 32'h42c64ce3, 32'hc2bc6526, 32'h428b1b4e, 32'hc231171b, 32'hc2716a3d, 32'h42649e5c, 32'h40728c7a};
test_label[4002] = '{32'h42649e5c};
test_output[4002] = '{32'h4227fb6b};
/*############ DEBUG ############
test_input[32016:32023] = '{75.1877111744, 99.1501713471, -94.1975583556, 69.5533257392, -44.272562901, -60.3537474016, 57.1546465249, 3.78982404804};
test_label[4002] = '{57.1546465249};
test_output[4002] = '{41.9955248222};
############ END DEBUG ############*/
test_input[32024:32031] = '{32'hc2775b4a, 32'hc145893a, 32'hc269f6e4, 32'hc292248d, 32'h42127049, 32'hc1e7a6ba, 32'h41260715, 32'hc25f9742};
test_label[4003] = '{32'h42127049};
test_output[4003] = '{32'h2c8e6900};
/*############ DEBUG ############
test_input[32024:32031] = '{-61.8391511366, -12.3460023486, -58.4911030001, -73.0713896375, 36.6096543613, -28.9564097244, 10.3767286067, -55.8977137666};
test_label[4003] = '{36.6096543613};
test_output[4003] = '{4.04754008088e-12};
############ END DEBUG ############*/
test_input[32032:32039] = '{32'h42990119, 32'h42c059e6, 32'hc2252259, 32'h42b98eef, 32'hc220ada2, 32'hc12e060d, 32'h3f2f705a, 32'hc18a2b43};
test_label[4004] = '{32'h42990119};
test_output[4004] = '{32'h419da6aa};
/*############ DEBUG ############
test_input[32032:32039] = '{76.5021469601, 96.1755816263, -41.283542672, 92.779163371, -40.1695649366, -10.8764776403, 0.685308074992, -17.2711230529};
test_label[4004] = '{76.5021469601};
test_output[4004] = '{19.7063790143};
############ END DEBUG ############*/
test_input[32040:32047] = '{32'hc13b880b, 32'hc095e5d8, 32'h42002bd8, 32'hc0d8ec0e, 32'h429b7598, 32'hc1b371eb, 32'h426ad975, 32'hc132e802};
test_label[4005] = '{32'h426ad975};
test_output[4005] = '{32'h41982378};
/*############ DEBUG ############
test_input[32040:32047] = '{-11.7207137835, -4.68430718103, 32.0428177323, -6.77881537173, 77.7296775142, -22.4306235092, 58.7123597205, -11.1816421435};
test_label[4005] = '{58.7123597205};
test_output[4005] = '{19.0173177992};
############ END DEBUG ############*/
test_input[32048:32055] = '{32'h41a43f50, 32'h42098906, 32'hc255e586, 32'hc2688eb7, 32'hc2887155, 32'h411010e9, 32'hc117efb4, 32'h429a5b39};
test_label[4006] = '{32'hc2688eb7};
test_output[4006] = '{32'h4307514a};
/*############ DEBUG ############
test_input[32048:32055] = '{20.530914502, 34.3838134613, -53.474142595, -58.1393695139, -68.2213493791, 9.00412831583, -9.49602125662, 77.1781668721};
test_label[4006] = '{-58.1393695139};
test_output[4006] = '{135.317536386};
############ END DEBUG ############*/
test_input[32056:32063] = '{32'h41f64360, 32'h42989c19, 32'hc23edbe5, 32'h42061016, 32'h42839347, 32'h42c0de71, 32'h41983adc, 32'hc285e45c};
test_label[4007] = '{32'h41983adc};
test_output[4007] = '{32'h429acfba};
/*############ DEBUG ############
test_input[32056:32063] = '{30.7828984432, 76.3048818437, -47.7147402991, 33.5157103919, 65.7876518517, 96.4344526934, 19.0287401574, -66.9460132851};
test_label[4007] = '{19.0287401574};
test_output[4007] = '{77.4057125378};
############ END DEBUG ############*/
test_input[32064:32071] = '{32'h416465e7, 32'hc293b2ae, 32'h41d4fb55, 32'h403eff89, 32'hc268155c, 32'hc28c07fd, 32'hc2380f59, 32'h4166c8bf};
test_label[4008] = '{32'h41d4fb55};
test_output[4008] = '{32'h371d4ddc};
/*############ DEBUG ############
test_input[32064:32071] = '{14.2748780263, -73.8489813913, 26.6227213161, 2.9843466155, -58.0208605276, -70.0156003617, -46.0149876386, 14.4240106332};
test_label[4008] = '{26.6227213161};
test_output[4008] = '{9.37605725074e-06};
############ END DEBUG ############*/
test_input[32072:32079] = '{32'hc2c7b898, 32'h41260b4f, 32'h42c3b778, 32'h41c60619, 32'h42967d78, 32'hc224199c, 32'h41f123b9, 32'hc1d04d14};
test_label[4009] = '{32'h41f123b9};
test_output[4009] = '{32'h42876e89};
/*############ DEBUG ############
test_input[32072:32079] = '{-99.8605326015, 10.3777605321, 97.8583345458, 24.7529778452, 75.24505434, -41.0250097688, 30.1424433252, -26.0376349036};
test_label[4009] = '{30.1424433252};
test_output[4009] = '{67.7158912208};
############ END DEBUG ############*/
test_input[32080:32087] = '{32'h4256c0ef, 32'h423d3c31, 32'h42b1d5e3, 32'h42670478, 32'h428aa202, 32'hc1f5a655, 32'h425434b7, 32'h41c2a2e7};
test_label[4010] = '{32'h4256c0ef};
test_output[4010] = '{32'h420cead7};
/*############ DEBUG ############
test_input[32080:32087] = '{53.688410118, 47.3087789813, 88.9177476425, 57.7543654552, 69.3164207934, -30.7062176207, 53.0514808867, 24.3295418988};
test_label[4010] = '{53.688410118};
test_output[4010] = '{35.2293375277};
############ END DEBUG ############*/
test_input[32088:32095] = '{32'h41d9ac63, 32'h42ab160d, 32'hc2b1f1f3, 32'hc296da93, 32'hc2b6b940, 32'h42bcc78d, 32'hc2c2384f, 32'h428ed7be};
test_label[4011] = '{32'h42bcc78d};
test_output[4011] = '{32'h3916d5d3};
/*############ DEBUG ############
test_input[32088:32095] = '{27.2091722739, 85.5430641935, -88.9725577465, -75.426900893, -91.3618149043, 94.3897484439, -97.1099742256, 71.4213719385};
test_label[4011] = '{94.3897484439};
test_output[4011] = '{0.000143847702599};
############ END DEBUG ############*/
test_input[32096:32103] = '{32'hc26b01f1, 32'h4124cb8a, 32'h414e2ffd, 32'h409732e2, 32'h42c6126c, 32'h42a3e6bc, 32'h425aea97, 32'hc288589a};
test_label[4012] = '{32'h409732e2};
test_output[4012] = '{32'h42bc9f3e};
/*############ DEBUG ############
test_input[32096:32103] = '{-58.7518965398, 10.2996923189, 12.8867159479, 4.7249611416, 99.0359778016, 81.9506532224, 54.7290924909, -68.1730530394};
test_label[4012] = '{4.7249611416};
test_output[4012] = '{94.311016698};
############ END DEBUG ############*/
test_input[32104:32111] = '{32'h42940547, 32'h4280854e, 32'h41a78bd0, 32'h42880b93, 32'hc290d153, 32'hc20f1db8, 32'h410cfd61, 32'h421bf5f4};
test_label[4013] = '{32'h42940547};
test_output[4013] = '{32'h3b28101b};
/*############ DEBUG ############
test_input[32104:32111] = '{74.0103061098, 64.2603591263, 20.9432679263, 68.0226063688, -72.4088383808, -35.7790216156, 8.81185982369, 38.9901876646};
test_label[4013] = '{74.0103061098};
test_output[4013] = '{0.00256443652925};
############ END DEBUG ############*/
test_input[32112:32119] = '{32'h4271ab85, 32'hc26766c7, 32'hc184d772, 32'hc151800b, 32'hc1a342a9, 32'h428bfd20, 32'h418ee4f6, 32'hc2bad64d};
test_label[4014] = '{32'hc184d772};
test_output[4014] = '{32'h42ad3305};
/*############ DEBUG ############
test_input[32112:32119] = '{60.4175003821, -57.8503695268, -16.6051977326, -13.0937604496, -20.4075489473, 69.9943827539, 17.8617965551, -93.4185545782};
test_label[4014] = '{-16.6051977326};
test_output[4014] = '{86.5996497968};
############ END DEBUG ############*/
test_input[32120:32127] = '{32'hc220e664, 32'hc2834241, 32'h424ba2c9, 32'h425c4553, 32'h4293a131, 32'h42a7ec3b, 32'h42613f34, 32'h42429636};
test_label[4015] = '{32'h42a7ec3b};
test_output[4015] = '{32'h38247571};
/*############ DEBUG ############
test_input[32120:32127] = '{-40.2249895921, -65.629405113, 50.9089707152, 55.0677005411, 73.8148255949, 83.9613841728, 56.3117228398, 48.6466905333};
test_label[4015] = '{83.9613841728};
test_output[4015] = '{3.92100231767e-05};
############ END DEBUG ############*/
test_input[32128:32135] = '{32'h41dfb7cc, 32'h428cc789, 32'h42bd038c, 32'hc2083550, 32'hc22e5da7, 32'hc2b281f7, 32'h424fb198, 32'h426cebe1};
test_label[4016] = '{32'h41dfb7cc};
test_output[4016] = '{32'h42851599};
/*############ DEBUG ############
test_input[32128:32135] = '{27.9647447531, 70.389718246, 94.5069272921, -34.052061088, -43.5914568464, -89.2538347108, 51.9234313188, 59.2303503321};
test_label[4016] = '{27.9647447531};
test_output[4016] = '{66.542182539};
############ END DEBUG ############*/
test_input[32136:32143] = '{32'hc227aa53, 32'hc21ee9c9, 32'h4210b881, 32'hc22e8bf7, 32'h42bc2bfd, 32'hc29787ec, 32'h4289000d, 32'h42ada3f2};
test_label[4017] = '{32'hc227aa53};
test_output[4017] = '{32'h430800c1};
/*############ DEBUG ############
test_input[32136:32143] = '{-41.9163324654, -39.7283065185, 36.1801800919, -43.6366847598, 94.0859162289, -75.7654740151, 68.5000954021, 86.8202042196};
test_label[4017] = '{-41.9163324654};
test_output[4017] = '{136.002947553};
############ END DEBUG ############*/
test_input[32144:32151] = '{32'h40d41107, 32'hc2aaa834, 32'hc1e7c343, 32'hc2c12305, 32'hc28e93d7, 32'hc2c5d2cb, 32'hc21caa7f, 32'h4287ea16};
test_label[4018] = '{32'hc28e93d7};
test_output[4018] = '{32'h430b3ef7};
/*############ DEBUG ############
test_input[32144:32151] = '{6.62707835994, -85.3285241385, -28.9703424158, -96.568394535, -71.2887532074, -98.9117040798, -39.166501623, 67.9572007745};
test_label[4018] = '{-71.2887532074};
test_output[4018] = '{139.245953982};
############ END DEBUG ############*/
test_input[32152:32159] = '{32'h4149c075, 32'hc162be80, 32'hc081d31c, 32'h417fa240, 32'h4224abab, 32'hc2259ee6, 32'h42b15bb0, 32'h42b4dd74};
test_label[4019] = '{32'h42b15bb0};
test_output[4019] = '{32'h3ff4e27a};
/*############ DEBUG ############
test_input[32152:32159] = '{12.6094865806, -14.171508866, -4.05702032781, 15.9771115968, 41.1676441334, -41.4051733819, 88.6790793241, 90.4325262293};
test_label[4019] = '{88.6790793241};
test_output[4019] = '{1.91316149971};
############ END DEBUG ############*/
test_input[32160:32167] = '{32'h42671577, 32'hbfb3864b, 32'h42389c00, 32'h42953ed1, 32'h4262f39a, 32'hc171f684, 32'hc26a8c76, 32'h42bcd40b};
test_label[4020] = '{32'hbfb3864b};
test_output[4020] = '{32'h42bfa224};
/*############ DEBUG ############
test_input[32160:32167] = '{57.7709625282, -1.40253585435, 46.1523435408, 74.6226909545, 56.7378915953, -15.1226847602, -58.6371687656, 94.4141477614};
test_label[4020] = '{-1.40253585435};
test_output[4020] = '{95.8166836183};
############ END DEBUG ############*/
test_input[32168:32175] = '{32'h42bf8fb6, 32'hc14b4732, 32'hc20c0d3d, 32'h41e9fe78, 32'hc1866376, 32'h4287b60c, 32'hc10e9445, 32'h429221e5};
test_label[4021] = '{32'hc14b4732};
test_output[4021] = '{32'h42d8f89d};
/*############ DEBUG ############
test_input[32168:32175] = '{95.7806881673, -12.7048820284, -35.0129272736, 29.2492529498, -16.7985648985, 67.8555578676, -8.91119845171, 73.066203328};
test_label[4021] = '{-12.7048820284};
test_output[4021] = '{108.485570196};
############ END DEBUG ############*/
test_input[32176:32183] = '{32'hbf8ea232, 32'h428c0cff, 32'hc230cceb, 32'hc28c10d0, 32'hc2578f4a, 32'hc237ad33, 32'h42b576cb, 32'h42bbc1e0};
test_label[4022] = '{32'hc237ad33};
test_output[4022] = '{32'h430bd704};
/*############ DEBUG ############
test_input[32176:32183] = '{-1.11432483493, 70.0253813849, -44.2001159743, -70.0328372277, -53.88993172, -45.9191393539, 90.7320168817, 93.8786608712};
test_label[4022] = '{-45.9191393539};
test_output[4022] = '{139.839897739};
############ END DEBUG ############*/
test_input[32184:32191] = '{32'h42a38434, 32'h4282ff47, 32'h42c28252, 32'hc281379a, 32'h42579f09, 32'h41540a28, 32'hc2a2da91, 32'hc11c28d3};
test_label[4023] = '{32'hc281379a};
test_output[4023] = '{32'h4321dcf6};
/*############ DEBUG ############
test_input[32184:32191] = '{81.7582085772, 65.4985849618, 97.25453103, -64.6085962445, 53.9053061225, 13.252480016, -81.4268905941, -9.75996722895};
test_label[4023] = '{-64.6085962445};
test_output[4023] = '{161.863127461};
############ END DEBUG ############*/
test_input[32192:32199] = '{32'h41c122d9, 32'h4286061f, 32'h42829653, 32'h420b4e2a, 32'hc2acc5d6, 32'hc1bb6946, 32'h41e276da, 32'h421b0b6a};
test_label[4024] = '{32'h41c122d9};
test_output[4024] = '{32'h422c23c1};
/*############ DEBUG ############
test_input[32192:32199] = '{24.1420161534, 67.0119588732, 65.2936008182, 34.8263331389, -86.386396407, -23.4264033355, 28.3080327971, 38.7611453549};
test_label[4024] = '{24.1420161534};
test_output[4024] = '{43.0349149827};
############ END DEBUG ############*/
test_input[32200:32207] = '{32'hbea8a5f3, 32'h428a7088, 32'hc2abbaf3, 32'h41fa17ec, 32'h410fd5f4, 32'hc1c1bdf7, 32'hc2c4f354, 32'h4276cf21};
test_label[4025] = '{32'h4276cf21};
test_output[4025] = '{32'h40f093ed};
/*############ DEBUG ############
test_input[32200:32207] = '{-0.329391096873, 69.21978837, -85.8651365697, 31.2616813595, 8.98973433193, -24.2177555113, -98.4752469487, 61.7022742503};
test_label[4025] = '{61.7022742503};
test_output[4025] = '{7.51805745403};
############ END DEBUG ############*/
test_input[32208:32215] = '{32'h428cc1b4, 32'hc1b2e850, 32'h420667fa, 32'h418ffddb, 32'h426c3ae0, 32'hc2a450fe, 32'h4297371e, 32'h42570552};
test_label[4026] = '{32'hc2a450fe};
test_output[4026] = '{32'h431dc56c};
/*############ DEBUG ############
test_input[32208:32215] = '{70.3783258689, -22.3634339981, 33.601540233, 17.9989536945, 59.0574936248, -82.1581886693, 75.6076530406, 53.7551949613};
test_label[4026] = '{-82.1581886693};
test_output[4026] = '{157.771184605};
############ END DEBUG ############*/
test_input[32216:32223] = '{32'hc220b455, 32'hc23433a7, 32'h42b0632c, 32'hc26801be, 32'h42692ed7, 32'h420d7122, 32'hc28883f5, 32'h420a4c43};
test_label[4027] = '{32'hc23433a7};
test_output[4027] = '{32'h43053e80};
/*############ DEBUG ############
test_input[32216:32223] = '{-40.1761055101, -45.0504432025, 88.193695329, -58.0017022306, 58.2957419626, 35.3604799678, -68.2577248494, 34.5744740025};
test_label[4027] = '{-45.0504432025};
test_output[4027] = '{133.244138531};
############ END DEBUG ############*/
test_input[32224:32231] = '{32'hc1ddfa90, 32'h426c75b1, 32'hc26f4283, 32'hc234f4c5, 32'h42a0af15, 32'hc1888575, 32'hc2470c3c, 32'h42a21239};
test_label[4028] = '{32'hc1ddfa90};
test_output[4028] = '{32'h42da6060};
/*############ DEBUG ############
test_input[32224:32231] = '{-27.7473446119, 59.114933258, -59.8149541949, -45.2390314118, 80.3419537952, -17.0651640129, -49.7619470833, 81.0355891733};
test_label[4028] = '{-27.7473446119};
test_output[4028] = '{109.188236188};
############ END DEBUG ############*/
test_input[32232:32239] = '{32'hc27e2614, 32'hc13940c2, 32'h4213745f, 32'hc2b29685, 32'hc2699703, 32'h42aa1e85, 32'hc1ec4c5a, 32'h422b10db};
test_label[4029] = '{32'h42aa1e85};
test_output[4029] = '{32'h80000000};
/*############ DEBUG ############
test_input[32232:32239] = '{-63.5371874933, -11.5783103658, 36.8636451834, -89.2939834527, -58.3974715755, 85.0596049122, -29.5372810407, 42.7664620951};
test_label[4029] = '{85.0596049122};
test_output[4029] = '{-0.0};
############ END DEBUG ############*/
test_input[32240:32247] = '{32'hc26fcafa, 32'hc299dcab, 32'hc2b7d83a, 32'h428681f2, 32'h41d7c686, 32'hc2acdfb0, 32'hc2893e8f, 32'hc29e9f04};
test_label[4030] = '{32'hc2893e8f};
test_output[4030] = '{32'h4307e041};
/*############ DEBUG ############
test_input[32240:32247] = '{-59.9482187816, -76.930994448, -91.9223168015, 67.2538016458, 26.9719357367, -86.4368866026, -68.6221839897, -79.3105772782};
test_label[4030] = '{-68.6221839897};
test_output[4030] = '{135.875985635};
############ END DEBUG ############*/
test_input[32248:32255] = '{32'hc19a687f, 32'hc2c24b12, 32'h41fe4aa4, 32'hc2b4239e, 32'hc2af006a, 32'h41dd8ef2, 32'h40190673, 32'h41bf546c};
test_label[4031] = '{32'hc2b4239e};
test_output[4031] = '{32'h42f3bef5};
/*############ DEBUG ############
test_input[32248:32255] = '{-19.3010230331, -97.1466247871, 31.7864449742, -90.0695653166, -87.5008114539, 27.6947981716, 2.39101861239, 23.9162218114};
test_label[4031] = '{-90.0695653166};
test_output[4031] = '{121.872959478};
############ END DEBUG ############*/
test_input[32256:32263] = '{32'hc23be3b9, 32'h409e69a1, 32'hc013fc3c, 32'h4229fb30, 32'h41b4eb88, 32'hbfaa00d5, 32'h41d3776c, 32'h4048b9f7};
test_label[4032] = '{32'h4048b9f7};
test_output[4032] = '{32'h421d6f90};
/*############ DEBUG ############
test_input[32256:32263] = '{-46.9723857913, 4.9503940637, -2.31227018747, 42.4952985798, 22.6150057693, -1.32815035472, 26.433312176, 3.13635050302};
test_label[4032] = '{3.13635050302};
test_output[4032] = '{39.3589481849};
############ END DEBUG ############*/
test_input[32264:32271] = '{32'hc009e714, 32'hc2985cdd, 32'h42898d53, 32'hc2bba7df, 32'hc1406c2b, 32'hc2286ac9, 32'hc2a68f8c, 32'hc2740dfc};
test_label[4033] = '{32'hc2985cdd};
test_output[4033] = '{32'h4310f518};
/*############ DEBUG ############
test_input[32264:32271] = '{-2.15472891434, -76.181374048, 68.7760229528, -93.8278718926, -12.026407808, -42.1042822693, -83.2803637883, -61.0136564634};
test_label[4033] = '{-76.181374048};
test_output[4033] = '{144.957397001};
############ END DEBUG ############*/
test_input[32272:32279] = '{32'h41ec3b7a, 32'h42a1a8ee, 32'hc238ec58, 32'hc2acc7da, 32'hc082a3da, 32'hc2c7955f, 32'h42816e17, 32'hc2ab10f6};
test_label[4034] = '{32'hc082a3da};
test_output[4034] = '{32'h42a9d32c};
/*############ DEBUG ############
test_input[32272:32279] = '{29.529040677, 80.8299416715, -46.2308035335, -86.3903320551, -4.08250139146, -99.7917384078, 64.7150226668, -85.5331292597};
test_label[4034] = '{-4.08250139146};
test_output[4034] = '{84.9124431633};
############ END DEBUG ############*/
test_input[32280:32287] = '{32'h42ac5496, 32'hc26c987c, 32'h429f7583, 32'h405ce357, 32'hc2846461, 32'hc2b361e3, 32'hc1e9adca, 32'h425ad2d2};
test_label[4035] = '{32'hc2846461};
test_output[4035] = '{32'h43185ce4};
/*############ DEBUG ############
test_input[32280:32287] = '{86.1652063826, -59.148908996, 79.7295187238, 3.45137566037, -66.1960500468, -89.6911832149, -29.2098570165, 54.7058808048};
test_label[4035] = '{-66.1960500468};
test_output[4035] = '{152.362858451};
############ END DEBUG ############*/
test_input[32288:32295] = '{32'h416dbd80, 32'hc28a9380, 32'hc204448c, 32'hc2b77cc0, 32'hc2abf668, 32'hc10dbb72, 32'h41c0a3c2, 32'h42c7e29e};
test_label[4036] = '{32'h416dbd80};
test_output[4036] = '{32'h42aa2aee};
/*############ DEBUG ############
test_input[32288:32295] = '{14.8587648814, -69.2880888897, -33.0669404071, -91.7436559062, -85.9812589712, -8.85826297902, 24.0799603148, 99.9426119855};
test_label[4036] = '{14.8587648814};
test_output[4036] = '{85.0838471041};
############ END DEBUG ############*/
test_input[32296:32303] = '{32'hc2c47726, 32'hc2a5ee8d, 32'hc263433d, 32'h424dbcef, 32'h40de1f38, 32'hc2562d97, 32'h41466288, 32'h429db52d};
test_label[4037] = '{32'h429db52d};
test_output[4037] = '{32'h2bade800};
/*############ DEBUG ############
test_input[32296:32303] = '{-98.2327083176, -82.9659171824, -56.815661889, 51.4345071656, 6.94131100071, -53.5445196451, 12.399055112, 78.8538619894};
test_label[4037] = '{78.8538619894};
test_output[4037] = '{1.23567822641e-12};
############ END DEBUG ############*/
test_input[32304:32311] = '{32'hc1b5932a, 32'h422d362e, 32'h422a3b57, 32'hc06651d8, 32'h42ab86d7, 32'h419f5101, 32'h42bbfa9b, 32'h42b430ef};
test_label[4038] = '{32'h42b430ef};
test_output[4038] = '{32'h407a8417};
/*############ DEBUG ############
test_input[32304:32311] = '{-22.6968572039, 43.3029102289, 42.5579499798, -3.59874526659, 85.7633577341, 19.9145526525, 93.9894627298, 90.0955741422};
test_label[4038] = '{90.0955741422};
test_output[4038] = '{3.91431217242};
############ END DEBUG ############*/
test_input[32312:32319] = '{32'h423a6619, 32'h427d1f6f, 32'h409727e9, 32'hc26a372c, 32'h429098cf, 32'h4290bbad, 32'hc280894b, 32'h4216e322};
test_label[4039] = '{32'h423a6619};
test_output[4039] = '{32'h41d369a5};
/*############ DEBUG ############
test_input[32312:32319] = '{46.5997039682, 63.280695314, 4.72362201098, -58.5538774143, 72.298454834, 72.3665515239, -64.2681502275, 37.7218079001};
test_label[4039] = '{46.5997039682};
test_output[4039] = '{26.4265844781};
############ END DEBUG ############*/
test_input[32320:32327] = '{32'hc29d39ac, 32'h4180fc28, 32'h42afe27f, 32'hc18b2f82, 32'h42854b10, 32'hc253aff4, 32'hc29bd59f, 32'h427ae620};
test_label[4040] = '{32'hc18b2f82};
test_output[4040] = '{32'h42d2ae5f};
/*############ DEBUG ############
test_input[32320:32327] = '{-78.6126403837, 16.1231228666, 87.9423758648, -17.3981962955, 66.6466099975, -52.9218304938, -77.9172314743, 62.7247316252};
test_label[4040] = '{-17.3981962955};
test_output[4040] = '{105.340572161};
############ END DEBUG ############*/
test_input[32328:32335] = '{32'hc2074366, 32'hc29ff97e, 32'h414b61b2, 32'h42bb8932, 32'hc246c1aa, 32'h42c34614, 32'hc2b918f8, 32'h3e8dadee};
test_label[4041] = '{32'hc29ff97e};
test_output[4041] = '{32'h4331a514};
/*############ DEBUG ############
test_input[32328:32335] = '{-33.8158187368, -79.9872899295, 12.7113515137, 93.7679610362, -49.689125762, 97.6368731363, -92.5487700583, 0.276717600751};
test_label[4041] = '{-79.9872899295};
test_output[4041] = '{177.644829118};
############ END DEBUG ############*/
test_input[32336:32343] = '{32'hc285208e, 32'h421f69ad, 32'h42aa3da2, 32'h42c1833c, 32'hc1a66379, 32'hc24151fd, 32'h40bc3266, 32'h418e950f};
test_label[4042] = '{32'h418e950f};
test_output[4042] = '{32'h429dddfa};
/*############ DEBUG ############
test_input[32336:32343] = '{-66.5635840778, 39.8531992287, 85.120376892, 96.7563193757, -20.7985712405, -48.330067883, 5.88115214782, 17.8227822816};
test_label[4042] = '{17.8227822816};
test_output[4042] = '{78.9335459366};
############ END DEBUG ############*/
test_input[32344:32351] = '{32'h424ef783, 32'h420c4cba, 32'hc11d8f85, 32'hc1893c42, 32'h41fa7e09, 32'hbf413d71, 32'h41cac6b8, 32'h421eb23a};
test_label[4043] = '{32'hbf413d71};
test_output[4043] = '{32'h4251fc7b};
/*############ DEBUG ############
test_input[32344:32351] = '{51.7417121763, 35.0749264743, -9.84753918679, -17.1544223558, 31.3115407523, -0.754843768113, 25.3470311503, 39.674048948};
test_label[4043] = '{-0.754843768113};
test_output[4043] = '{52.4965617457};
############ END DEBUG ############*/
test_input[32352:32359] = '{32'h428bebc3, 32'hc22bb0d7, 32'hc2bf6edb, 32'h417ee4f4, 32'h4120fb68, 32'h41ff3bd9, 32'h41ff3c8d, 32'hc18a1674};
test_label[4044] = '{32'hc2bf6edb};
test_output[4044] = '{32'h4325ad4f};
/*############ DEBUG ############
test_input[32352:32359] = '{69.9604751571, -42.9226946681, -95.7165157662, 15.9308966673, 10.0613780027, 31.9042234237, 31.9045653403, -17.260963102};
test_label[4044] = '{-95.7165157662};
test_output[4044] = '{165.676990923};
############ END DEBUG ############*/
test_input[32360:32367] = '{32'hc11b5aab, 32'h4240db8c, 32'hc2864b4e, 32'h42c04103, 32'hc20512bf, 32'hc00bdda3, 32'hc19b5914, 32'hc1de85f1};
test_label[4045] = '{32'hc11b5aab};
test_output[4045] = '{32'h42d3ac59};
/*############ DEBUG ############
test_input[32360:32367] = '{-9.7096356218, 48.2144003797, -67.1470830385, 96.1269784779, -33.2683068968, -2.18540263652, -19.4184945742, -27.8154003673};
test_label[4045] = '{-9.7096356218};
test_output[4045] = '{105.8366141};
############ END DEBUG ############*/
test_input[32368:32375] = '{32'h42aebb5a, 32'hc2aed273, 32'h41fdc079, 32'hc2c52d08, 32'h42394352, 32'h4227e891, 32'h428e3669, 32'h415cccd8};
test_label[4046] = '{32'hc2c52d08};
test_output[4046] = '{32'h4339f431};
/*############ DEBUG ############
test_input[32368:32375] = '{87.3659246104, -87.4110308734, 31.7189815875, -98.5879491892, 46.3157424022, 41.9771160241, 71.106273241, 13.800010596};
test_label[4046] = '{-98.5879491892};
test_output[4046] = '{185.953873886};
############ END DEBUG ############*/
test_input[32376:32383] = '{32'hc24b8e42, 32'h42a6b991, 32'h42943a3a, 32'h40bbb19b, 32'hc21bcd94, 32'h42c583b6, 32'h41f41418, 32'hc21db9ba};
test_label[4047] = '{32'h42943a3a};
test_output[4047] = '{32'h41c525ef};
/*############ DEBUG ############
test_input[32376:32383] = '{-50.8889235599, 83.3624319643, 74.1137250783, 5.86543051952, -38.9507606071, 98.7572475374, 30.5098117347, -39.4313738083};
test_label[4047] = '{74.1137250783};
test_output[4047] = '{24.6435226653};
############ END DEBUG ############*/
test_input[32384:32391] = '{32'h42c399a1, 32'h424f61a5, 32'hc21bf8e5, 32'hc203ae15, 32'hc1558f77, 32'hc12cc62e, 32'hc21b7639, 32'hc112d9aa};
test_label[4048] = '{32'hc112d9aa};
test_output[4048] = '{32'h42d5f4d7};
/*############ DEBUG ############
test_input[32384:32391] = '{97.8000587351, 51.8453549841, -38.9930601275, -32.9200025827, -13.3475259221, -10.798383361, -38.8654529798, -9.17814064232};
test_label[4048] = '{-9.17814064232};
test_output[4048] = '{106.978199377};
############ END DEBUG ############*/
test_input[32392:32399] = '{32'h4226f3a0, 32'hc17ce26b, 32'h4204786c, 32'hc1d79a87, 32'hc2b4ee02, 32'hc2864622, 32'h41714284, 32'h42b56890};
test_label[4049] = '{32'h4226f3a0};
test_output[4049] = '{32'h4243dd80};
/*############ DEBUG ############
test_input[32392:32399] = '{41.7379132476, -15.8052782661, 33.1175996231, -26.9504520851, -90.4648572338, -67.1369795092, 15.0787390957, 90.7042235554};
test_label[4049] = '{41.7379132476};
test_output[4049] = '{48.9663103078};
############ END DEBUG ############*/
test_input[32400:32407] = '{32'hc22543cb, 32'h409a1ab6, 32'hc208467d, 32'hc2ae7876, 32'hc0c8d7b8, 32'h420d0c1d, 32'h41af5d48, 32'hc24dbf41};
test_label[4050] = '{32'h420d0c1d};
test_output[4050] = '{32'h35d7a844};
/*############ DEBUG ############
test_input[32400:32407] = '{-41.3162041888, 4.81576048332, -34.0688349413, -87.2352761251, -6.27633288697, 35.2618302754, 21.9205476687, -51.436769739};
test_label[4050] = '{35.2618302754};
test_output[4050] = '{1.60677198047e-06};
############ END DEBUG ############*/
test_input[32408:32415] = '{32'h421b893d, 32'h4254704b, 32'h4104da6a, 32'h428d8839, 32'h42aa0aa5, 32'h40ab003f, 32'h421960c8, 32'hc1981124};
test_label[4051] = '{32'h421960c8};
test_output[4051] = '{32'h423ab484};
/*############ DEBUG ############
test_input[32408:32415] = '{38.8840228752, 53.1096607573, 8.30332375769, 70.7660591242, 85.0207937951, 5.34378002447, 38.34451139, -19.0083698741};
test_label[4051] = '{38.34451139};
test_output[4051] = '{46.6762830497};
############ END DEBUG ############*/
test_input[32416:32423] = '{32'hc2b2d292, 32'hc22a18f0, 32'hc2a424b5, 32'h42aa0de8, 32'h41b565c1, 32'hc24ce591, 32'h4255e407, 32'h4184ebb1};
test_label[4052] = '{32'hc2b2d292};
test_output[4052] = '{32'h432e703d};
/*############ DEBUG ############
test_input[32416:32423] = '{-89.4112673258, -42.5243520301, -82.071696135, 85.0271574797, 22.6746836545, -51.2241862636, 53.4726826932, 16.615083714};
test_label[4052] = '{-89.4112673258};
test_output[4052] = '{174.438424805};
############ END DEBUG ############*/
test_input[32424:32431] = '{32'h42118f37, 32'h42504617, 32'h41cfe77e, 32'h4007cd39, 32'h422eb150, 32'h4197b2bb, 32'h42898046, 32'h4248665b};
test_label[4053] = '{32'h42898046};
test_output[4053] = '{32'h338b4520};
/*############ DEBUG ############
test_input[32424:32431] = '{36.3898569924, 52.0684484189, 25.9880335794, 2.12190082323, 43.6731554763, 18.9622711746, 68.750530865, 50.0999546975};
test_label[4053] = '{68.750530865};
test_output[4053] = '{6.48526580151e-08};
############ END DEBUG ############*/
test_input[32432:32439] = '{32'h429b3dc1, 32'hc173cab6, 32'hc08f8551, 32'h423c7ebe, 32'hc241b048, 32'h41aae756, 32'hc26d1532, 32'h422d5144};
test_label[4054] = '{32'h429b3dc1};
test_output[4054] = '{32'h29830000};
/*############ DEBUG ############
test_input[32432:32439] = '{77.620613995, -15.2369898329, -4.48502393075, 47.1237710061, -48.4221503723, 21.3629570537, -59.2706999476, 43.3293623118};
test_label[4054] = '{77.620613995};
test_output[4054] = '{5.81756864904e-14};
############ END DEBUG ############*/
test_input[32440:32447] = '{32'hc245046c, 32'h41e16192, 32'hc2276dc1, 32'hc1b0997b, 32'hc28b5b1e, 32'hc191f71e, 32'h42ac6ce1, 32'h42a9657b};
test_label[4055] = '{32'hc245046c};
test_output[4055] = '{32'h4307aa70};
/*############ DEBUG ############
test_input[32440:32447] = '{-49.2543182449, 28.1726414388, -41.8571810758, -22.074941293, -69.6779664733, -18.2456621546, 86.2126560278, 84.6982075616};
test_label[4055] = '{-49.2543182449};
test_output[4055] = '{135.665767302};
############ END DEBUG ############*/
test_input[32448:32455] = '{32'h40b6e780, 32'h4272f5b4, 32'hc29d639b, 32'hc2a12000, 32'hc2190fa6, 32'h42c024ae, 32'hc23ab526, 32'hc27294a4};
test_label[4056] = '{32'h4272f5b4};
test_output[4056] = '{32'h420d53a9};
/*############ DEBUG ############
test_input[32448:32455] = '{5.7157592251, 60.7399442244, -78.6945456386, -80.5624981046, -38.2652816445, 96.0716436866, -46.6769028207, -60.6451587239};
test_label[4056] = '{60.7399442244};
test_output[4056] = '{35.3316994622};
############ END DEBUG ############*/
test_input[32456:32463] = '{32'hbf16dd9e, 32'h425320cf, 32'hc21929b6, 32'hc29b3a69, 32'hc2bda2ab, 32'hc29a43a8, 32'hc24971da, 32'hc2a84510};
test_label[4057] = '{32'h425320cf};
test_output[4057] = '{32'h80000000};
/*############ DEBUG ############
test_input[32456:32463] = '{-0.589319088392, 52.782038931, -38.2907326522, -77.6140821221, -94.8177079069, -77.1321373869, -50.3611833102, -84.1348861264};
test_label[4057] = '{52.782038931};
test_output[4057] = '{-0.0};
############ END DEBUG ############*/
test_input[32464:32471] = '{32'hc26e4ede, 32'h411799a2, 32'hbfe227ac, 32'hc249c87e, 32'hc26cf997, 32'h420a3b8a, 32'h4202827d, 32'hbe3c206a};
test_label[4058] = '{32'hbfe227ac};
test_output[4058] = '{32'h4211d779};
/*############ DEBUG ############
test_input[32464:32471] = '{-59.5770200331, 9.4750081188, -1.76683567239, -50.4457922642, -59.2437395994, 34.5581453828, 32.627428146, -0.183717396131};
test_label[4058] = '{-1.76683567239};
test_output[4058] = '{36.4604242331};
############ END DEBUG ############*/
test_input[32472:32479] = '{32'h4298f2d5, 32'hc2860b3a, 32'h41aea27a, 32'hc28bab95, 32'h42255861, 32'hc22b19e8, 32'h42635e95, 32'hc22e1ffa};
test_label[4059] = '{32'h42255861};
test_output[4059] = '{32'h420c8d4a};
/*############ DEBUG ############
test_input[32472:32479] = '{76.4742842373, -67.0219235605, 21.829333463, -69.8351211638, 41.3363074285, -42.7752998019, 56.8423653298, -43.5312273857};
test_label[4059] = '{41.3363074285};
test_output[4059] = '{35.1379768118};
############ END DEBUG ############*/
test_input[32480:32487] = '{32'hc2a139c7, 32'hc09b900f, 32'h418aa1b5, 32'h4268514b, 32'h42afd1c2, 32'hbfc4249a, 32'hc2a35bc5, 32'hc2b38cef};
test_label[4060] = '{32'hbfc4249a};
test_output[4060] = '{32'h42b2e254};
/*############ DEBUG ############
test_input[32480:32487] = '{-80.6128499186, -4.86133548426, 17.3289594532, 58.0793869841, 87.9096814109, -1.53236704387, -81.6792407608, -89.7752615366};
test_label[4060] = '{-1.53236704387};
test_output[4060] = '{89.4420484548};
############ END DEBUG ############*/
test_input[32488:32495] = '{32'h3f8eadd6, 32'hc29749f6, 32'h41224d69, 32'hc28d250c, 32'h428c8f06, 32'hc2c5bbab, 32'hc22149e9, 32'h41d14b4a};
test_label[4061] = '{32'h41d14b4a};
test_output[4061] = '{32'h42307867};
/*############ DEBUG ############
test_input[32488:32495] = '{1.1146800452, -75.6444536284, 10.1438985168, -70.5723572025, 70.2793432815, -98.8665399889, -40.322178739, 26.1617629061};
test_label[4061] = '{26.1617629061};
test_output[4061] = '{44.1175803754};
############ END DEBUG ############*/
test_input[32496:32503] = '{32'hc2110864, 32'h41255a99, 32'h427c0a89, 32'hc192c868, 32'h41aaf627, 32'hc251a9e1, 32'hc21022b8, 32'hc0edfbea};
test_label[4062] = '{32'h427c0a89};
test_output[4062] = '{32'h80000000};
/*############ DEBUG ############
test_input[32496:32503] = '{-36.2581944859, 10.3346186441, 63.010289371, -18.3478537403, 21.3701920931, -52.4158964658, -36.0339045717, -7.43700126477};
test_label[4062] = '{63.010289371};
test_output[4062] = '{-0.0};
############ END DEBUG ############*/
test_input[32504:32511] = '{32'h42ae480c, 32'hc1e553a7, 32'hc233a22f, 32'hc2a657c9, 32'h421653c9, 32'h415245b1, 32'hc24a782c, 32'h4202353b};
test_label[4063] = '{32'hc2a657c9};
test_output[4063] = '{32'h432a4fea};
/*############ DEBUG ############
test_input[32504:32511] = '{87.1407132402, -28.6658464186, -44.9083815307, -83.1714571233, 37.581820624, 13.142014849, -50.6173553237, 32.551983881};
test_label[4063] = '{-83.1714571233};
test_output[4063] = '{170.312170364};
############ END DEBUG ############*/
test_input[32512:32519] = '{32'hc21df8b9, 32'h3f502a50, 32'hc1bc7ca0, 32'h4194bd83, 32'h42a11802, 32'h428e7bb1, 32'h429b1c97, 32'hc29896d9};
test_label[4064] = '{32'hc1bc7ca0};
test_output[4064] = '{32'h42d0504d};
/*############ DEBUG ############
test_input[32512:32519] = '{-39.492893097, 0.813145646249, -23.560852581, 18.5925348523, 80.5468875837, 71.2415862052, 77.5558389647, -76.2946256917};
test_label[4064] = '{-23.560852581};
test_output[4064] = '{104.156840445};
############ END DEBUG ############*/
test_input[32520:32527] = '{32'h41a0876f, 32'h422896b9, 32'h42401462, 32'h4163ae89, 32'h42c25cf0, 32'h4203f5cf, 32'hc0048c9f, 32'hc2aff87b};
test_label[4065] = '{32'h41a0876f};
test_output[4065] = '{32'h429a3b14};
/*############ DEBUG ############
test_input[32520:32527] = '{20.0661297266, 42.1471891931, 48.0199062244, 14.2301113295, 97.1815194502, 32.9900464553, -2.07108271847, -87.9853111358};
test_label[4065] = '{20.0661297266};
test_output[4065] = '{77.1153897236};
############ END DEBUG ############*/
test_input[32528:32535] = '{32'h428e00e3, 32'hc2171e35, 32'h42a887fc, 32'h42b20b63, 32'hc2b1b629, 32'h4227641c, 32'h428c37ed, 32'hc248c6bd};
test_label[4066] = '{32'hc2171e35};
test_output[4066] = '{32'h42fd9edf};
/*############ DEBUG ############
test_input[32528:32535] = '{71.001730995, -37.7794971771, 84.2655957666, 89.0222402476, -88.8557819255, 41.8477645222, 70.1092320826, -50.1940786519};
test_label[4066] = '{-37.7794971771};
test_output[4066] = '{126.810295124};
############ END DEBUG ############*/
test_input[32536:32543] = '{32'h41ae4aa3, 32'h42329db2, 32'h4247d75e, 32'h4288031a, 32'hc13f06ea, 32'hc2975180, 32'h426e1ae0, 32'h429ade0c};
test_label[4067] = '{32'h4288031a};
test_output[4067] = '{32'h4116d7e9};
/*############ DEBUG ############
test_input[32536:32543] = '{21.7864438063, 44.6540004724, 49.9603203005, 68.0060556868, -11.9391879572, -75.6591815376, 59.5262450631, 77.4336877576};
test_label[4067] = '{68.0060556868};
test_output[4067] = '{9.42771255384};
############ END DEBUG ############*/
test_input[32544:32551] = '{32'h42182cee, 32'hc104d056, 32'hc2bf95a1, 32'hc2850d97, 32'hc24fcbb9, 32'h40199f55, 32'h4299b849, 32'h42a1bfab};
test_label[4068] = '{32'hc2850d97};
test_output[4068] = '{32'h43136b35};
/*############ DEBUG ############
test_input[32544:32551] = '{38.0438782498, -8.30086285646, -95.7922461716, -66.5265415171, -51.9489493572, 2.40034983236, 76.8599351198, 80.8743509224};
test_label[4068] = '{-66.5265415171};
test_output[4068] = '{147.418784909};
############ END DEBUG ############*/
test_input[32552:32559] = '{32'hc2c440c9, 32'h402fda9a, 32'hc2b6006a, 32'hc2a3047d, 32'hc2070818, 32'h42629982, 32'h42c2487d, 32'hc2bd3114};
test_label[4069] = '{32'h402fda9a};
test_output[4069] = '{32'h42bcc9a8};
/*############ DEBUG ############
test_input[32552:32559] = '{-98.1265333133, 2.74771741651, -91.0008088211, -81.5087692834, -33.7579039088, 56.6499085247, 97.1415786204, -94.5958557388};
test_label[4069] = '{2.74771741651};
test_output[4069] = '{94.3938612038};
############ END DEBUG ############*/
test_input[32560:32567] = '{32'hc139ab03, 32'h4111b19e, 32'hc27a68cb, 32'hc2a82d57, 32'h42b1c2e4, 32'h42576c9c, 32'hc26d87c8, 32'h427e11ae};
test_label[4070] = '{32'hc2a82d57};
test_output[4070] = '{32'h432cf81e};
/*############ DEBUG ############
test_input[32560:32567] = '{-11.6042508253, 9.10586319131, -62.6023376637, -84.0885530678, 88.8806486266, 53.8560647657, -59.3825980155, 63.5172660284};
test_label[4070] = '{-84.0885530678};
test_output[4070] = '{172.969201694};
############ END DEBUG ############*/
test_input[32568:32575] = '{32'hc2af29eb, 32'h427b8aa1, 32'h42a6619c, 32'hc273db10, 32'h4136d31f, 32'h414afb81, 32'h4296fcff, 32'h4248341b};
test_label[4071] = '{32'hc273db10};
test_output[4071] = '{32'h431027b0};
/*############ DEBUG ############
test_input[32568:32575] = '{-87.5818690364, 62.8853793517, 83.1906417276, -60.9639275731, 11.4265432189, 12.6864021087, 75.494131393, 50.0508850832};
test_label[4071] = '{-60.9639275731};
test_output[4071] = '{144.155023609};
############ END DEBUG ############*/
test_input[32576:32583] = '{32'h42991a3a, 32'hc2c40967, 32'hc295dc86, 32'h42886cdb, 32'h4220e226, 32'hc22325d6, 32'h41bd0513, 32'h4225909f};
test_label[4072] = '{32'h4225909f};
test_output[4072] = '{32'h420ca414};
/*############ DEBUG ############
test_input[32576:32583] = '{76.5512241978, -98.0183636861, -74.9307109782, 68.2126086229, 40.220849596, -40.7869491929, 23.6274772178, 41.391232141};
test_label[4072] = '{41.391232141};
test_output[4072] = '{35.1602311314};
############ END DEBUG ############*/
test_input[32584:32591] = '{32'h425df15e, 32'hc28ecebc, 32'hc2c63b11, 32'hc281ca12, 32'h42a3f78f, 32'h41d76e92, 32'h425c16e1, 32'hc2a74359};
test_label[4073] = '{32'hc28ecebc};
test_output[4073] = '{32'h43196326};
/*############ DEBUG ############
test_input[32584:32591] = '{55.4857098753, -71.4037803198, -99.1153621007, -64.8946655441, 81.9835107843, 26.9289891558, 55.0223445343, -83.6315364783};
test_label[4073] = '{-71.4037803198};
test_output[4073] = '{153.387291104};
############ END DEBUG ############*/
test_input[32592:32599] = '{32'hc1083f23, 32'h42a9ffce, 32'hc2be375d, 32'hc24a1859, 32'h427e602a, 32'hc19dd412, 32'h4281b537, 32'h42bd4a11};
test_label[4074] = '{32'h42bd4a11};
test_output[4074] = '{32'h3887c6ef};
/*############ DEBUG ############
test_input[32592:32599] = '{-8.51541422669, 84.9996161593, -95.1081283106, -50.5237756303, 63.5939107685, -19.7285499757, 64.8539330683, 94.644660168};
test_label[4074] = '{94.644660168};
test_output[4074] = '{6.47435563345e-05};
############ END DEBUG ############*/
test_input[32600:32607] = '{32'h42a53c6c, 32'hc21b27d3, 32'h3ebdb2fd, 32'hc291b364, 32'h42a1ad49, 32'hc1200a8b, 32'hc24c5c5b, 32'h4105ef4e};
test_label[4075] = '{32'h3ebdb2fd};
test_output[4075] = '{32'h42a4ce8b};
/*############ DEBUG ############
test_input[32600:32607] = '{82.6180079051, -38.7888914111, 0.370506210107, -72.8503716499, 80.8384488933, -10.0025736571, -51.0901902275, 8.37092404481};
test_label[4075] = '{0.370506210107};
test_output[4075] = '{82.4034044371};
############ END DEBUG ############*/
test_input[32608:32615] = '{32'h4233a24d, 32'hc20f2b52, 32'h41b4af6a, 32'h42189566, 32'hc23ddc3b, 32'hc1ceed25, 32'hc2a24ee3, 32'h4291c8e5};
test_label[4076] = '{32'h4233a24d};
test_output[4076] = '{32'h41dfdefb};
/*############ DEBUG ############
test_input[32608:32615] = '{44.908497243, -35.792306416, 22.585651949, 38.1458952519, -47.4650698803, -25.8657930823, -81.1540764804, 72.8923744465};
test_label[4076] = '{44.908497243};
test_output[4076] = '{27.9838772035};
############ END DEBUG ############*/
test_input[32616:32623] = '{32'h4267d2a5, 32'hc21d748c, 32'h41de0cc4, 32'hc2adfbfa, 32'h42c2e78c, 32'hc26d6141, 32'h42511383, 32'h42ac8ea1};
test_label[4077] = '{32'h42ac8ea1};
test_output[4077] = '{32'h4132c760};
/*############ DEBUG ############
test_input[32616:32623] = '{57.9557056852, -39.3638158952, 27.7562329664, -86.9921441208, 97.4522362413, -59.3449744855, 52.2690534273, 86.2785744321};
test_label[4077] = '{86.2785744321};
test_output[4077] = '{11.1736758482};
############ END DEBUG ############*/
test_input[32624:32631] = '{32'h42b5d7d8, 32'h42a128f1, 32'h409d1bef, 32'h41d39498, 32'hc2bdb53a, 32'hc2acaae9, 32'h42bf9a0f, 32'hc11d446c};
test_label[4078] = '{32'hc2bdb53a};
test_output[4078] = '{32'h433ea995};
/*############ DEBUG ############
test_input[32624:32631] = '{90.9215720797, 80.5799607681, 4.9096599858, 26.4475553951, -94.8539611328, -86.3338098289, 95.8008966053, -9.82920464087};
test_label[4078] = '{-94.8539611328};
test_output[4078] = '{190.662431378};
############ END DEBUG ############*/
test_input[32632:32639] = '{32'h429c01e3, 32'h425303e2, 32'hc2754f84, 32'h40b94015, 32'hc2269ed3, 32'hc1f89cd3, 32'h423851f6, 32'h42b435cc};
test_label[4079] = '{32'hc2754f84};
test_output[4079] = '{32'h43176ec7};
/*############ DEBUG ############
test_input[32632:32639] = '{78.0036886921, 52.7537921995, -61.3276508567, 5.78907265329, -41.6551002064, -31.0765734505, 46.0800418239, 90.1050698501};
test_label[4079] = '{-61.3276508567};
test_output[4079] = '{151.432726259};
############ END DEBUG ############*/
test_input[32640:32647] = '{32'hc2ba67a6, 32'h42a3febf, 32'hc1490759, 32'hbd1264d2, 32'h42507863, 32'h4262d92e, 32'hc2098ea4, 32'h4214bdae};
test_label[4080] = '{32'h42507863};
test_output[4080] = '{32'h41ef0a35};
/*############ DEBUG ############
test_input[32640:32647] = '{-93.2024393455, 81.9975498192, -12.5642940544, -0.0357406808605, 52.117565647, 56.7120879767, -34.3892985057, 37.1852349106};
test_label[4080] = '{52.117565647};
test_output[4080] = '{29.8799841722};
############ END DEBUG ############*/
test_input[32648:32655] = '{32'hc1086c2f, 32'hc2bed7e8, 32'h4196ff1d, 32'hc0a3a949, 32'h428471da, 32'h40e34817, 32'h41c8c4be, 32'hc2217839};
test_label[4081] = '{32'hc2bed7e8};
test_output[4081] = '{32'h4321a4e1};
/*############ DEBUG ############
test_input[32648:32655] = '{-8.52641218582, -95.4216950958, 18.8745661464, -5.11441462307, 66.2223698939, 7.10255005585, 25.096066321, -40.3674032839};
test_label[4081] = '{-95.4216950958};
test_output[4081] = '{161.64406499};
############ END DEBUG ############*/
test_input[32656:32663] = '{32'hc1a30e2f, 32'hc26a859f, 32'h423013ff, 32'hc260badf, 32'hc28b7c02, 32'h410920eb, 32'h42633bd6, 32'hc287e973};
test_label[4082] = '{32'hc1a30e2f};
test_output[4082] = '{32'h429a6177};
/*############ DEBUG ############
test_input[32656:32663] = '{-20.3819261685, -58.6304903018, 44.0195282193, -56.1824895089, -69.7422008023, 8.57053652147, 56.8084341421, -67.9559534205};
test_label[4082] = '{-20.3819261685};
test_output[4082] = '{77.1903631021};
############ END DEBUG ############*/
test_input[32664:32671] = '{32'hc16b0b05, 32'h422825b1, 32'h429262e9, 32'hc1c03423, 32'hc23ae94e, 32'h4203cf7c, 32'h4120d7d0, 32'hc26e391d};
test_label[4083] = '{32'hc16b0b05};
test_output[4083] = '{32'h42afc449};
/*############ DEBUG ############
test_input[32664:32671] = '{-14.6901899813, 42.0368076344, 73.1931816911, -24.0254566897, -46.7278351114, 32.9526232512, 10.0526885741, -59.5557739686};
test_label[4083] = '{-14.6901899813};
test_output[4083] = '{87.8833716724};
############ END DEBUG ############*/
test_input[32672:32679] = '{32'h42a7ab41, 32'h42b38b26, 32'hc1b21a8d, 32'hc28dfaec, 32'hc2c65453, 32'hc0483ac7, 32'h4129af5b, 32'hc2972cfa};
test_label[4084] = '{32'h4129af5b};
test_output[4084] = '{32'h429e5694};
/*############ DEBUG ############
test_input[32672:32679] = '{83.8344801847, 89.7717757601, -22.2629634356, -70.9900788076, -99.1646992352, -3.12858753386, 10.6053116574, -75.5878459467};
test_label[4084] = '{10.6053116574};
test_output[4084] = '{79.1690997836};
############ END DEBUG ############*/
test_input[32680:32687] = '{32'h4213a146, 32'hc0630a68, 32'hc2743563, 32'h4287d288, 32'hc218a01f, 32'h41d4257b, 32'hc2b3d597, 32'hbeaf4435};
test_label[4085] = '{32'h4287d288};
test_output[4085] = '{32'h291a8000};
/*############ DEBUG ############
test_input[32680:32687] = '{36.9074921352, -3.54751025662, -61.0521364039, 67.9111905937, -38.1563665236, 26.518301386, -89.9171713796, -0.342317239356};
test_label[4085] = '{67.9111905937};
test_output[4085] = '{3.43058914609e-14};
############ END DEBUG ############*/
test_input[32688:32695] = '{32'hc1ef43b5, 32'h423d0ac8, 32'hc14d63cc, 32'hc2456f67, 32'h42aa8138, 32'h42056639, 32'hc25be4d3, 32'h4222210d};
test_label[4086] = '{32'h4222210d};
test_output[4086] = '{32'h4232e162};
/*############ DEBUG ############
test_input[32688:32695] = '{-29.9080603609, 47.2605280134, -12.8368649399, -49.3587910486, 85.2523785302, 33.3498280611, -54.9734629613, 40.5322776417};
test_label[4086] = '{40.5322776417};
test_output[4086] = '{44.7201008885};
############ END DEBUG ############*/
test_input[32696:32703] = '{32'h42b266ab, 32'hc2bc6a9f, 32'h42b9c6e3, 32'h42a5bccb, 32'hc285611a, 32'hc21709fb, 32'h41a9686b, 32'hc2378ae1};
test_label[4087] = '{32'hc21709fb};
test_output[4087] = '{32'h4302ac47};
/*############ DEBUG ############
test_input[32696:32703] = '{89.200524177, -94.2082437358, 92.8884535321, 82.8687368562, -66.689647843, -37.7597447723, 21.1759862403, -45.885622948};
test_label[4087] = '{-37.7597447723};
test_output[4087] = '{130.672957527};
############ END DEBUG ############*/
test_input[32704:32711] = '{32'h42910f72, 32'h42a67203, 32'h422c5e9b, 32'h419944de, 32'hc2949965, 32'h4202a278, 32'h428c4f78, 32'hc22e36d5};
test_label[4088] = '{32'h42910f72};
test_output[4088] = '{32'h412b14a2};
/*############ DEBUG ############
test_input[32704:32711] = '{72.5301656566, 83.2226781724, 43.0923895678, 19.1586269088, -74.2995969816, 32.6586597169, 70.1552161827, -43.5535479698};
test_label[4088] = '{72.5301656566};
test_output[4088] = '{10.6925373428};
############ END DEBUG ############*/
test_input[32712:32719] = '{32'hc2088663, 32'hc291f720, 32'hc1a11d9d, 32'hc2223d92, 32'hc21e6285, 32'hc1c0c285, 32'hc21d1352, 32'hc2a701e4};
test_label[4089] = '{32'hc1c0c285};
test_output[4089] = '{32'h407e5e04};
/*############ DEBUG ############
test_input[32712:32719] = '{-34.1312355105, -72.9826627846, -20.1394601555, -40.5601258316, -39.5962086483, -24.0949800144, -39.2688656557, -83.5036893615};
test_label[4089] = '{-24.0949800144};
test_output[4089] = '{3.97448837332};
############ END DEBUG ############*/
test_input[32720:32727] = '{32'hc18bdaf2, 32'hc2451700, 32'h421352fa, 32'h421a293c, 32'hc17ed3d1, 32'h428f18ba, 32'h42a3332a, 32'h40f90cd7};
test_label[4090] = '{32'h421352fa};
test_output[4090] = '{32'h42331365};
/*############ DEBUG ############
test_input[32720:32727] = '{-17.4819071289, -49.2724617272, 36.8310336306, 38.5402665078, -15.9267132609, 71.5482961733, 81.5999304185, 7.78281742117};
test_label[4090] = '{36.8310336306};
test_output[4090] = '{44.7689399022};
############ END DEBUG ############*/
test_input[32728:32735] = '{32'hc29b46c1, 32'h42c30497, 32'h423e8b81, 32'hc17ac788, 32'hc2a04ec8, 32'h407e0734, 32'hc25699e3, 32'hbfd0604d};
test_label[4091] = '{32'hc17ac788};
test_output[4091] = '{32'h42e25d88};
/*############ DEBUG ############
test_input[32728:32735] = '{-77.638187615, 97.5089615838, 47.6362336473, -15.6737134794, -80.1538732895, 3.9691896664, -53.6502792684, -1.6279389058};
test_label[4091] = '{-15.6737134794};
test_output[4091] = '{113.182675063};
############ END DEBUG ############*/
test_input[32736:32743] = '{32'hc2375614, 32'h42a9c108, 32'h42a3167a, 32'h421f0830, 32'hc25c7e8e, 32'h427ba48c, 32'hc1ee2ec1, 32'hc2c4b17d};
test_label[4092] = '{32'hc2c4b17d};
test_output[4092] = '{32'h4337423c};
/*############ DEBUG ############
test_input[32736:32743] = '{-45.8340625463, 84.8770132059, 81.5438957831, 39.7579974379, -55.1235889197, 62.9106888429, -29.7728285925, -98.3466595073};
test_label[4092] = '{-98.3466595073};
test_output[4092] = '{183.258732567};
############ END DEBUG ############*/
test_input[32744:32751] = '{32'h41a10de6, 32'h42476d24, 32'h41be209d, 32'hc2778b81, 32'h422b6491, 32'h40c5a165, 32'h4036e33e, 32'h42054bbe};
test_label[4093] = '{32'h41a10de6};
test_output[4093] = '{32'h41edce3b};
/*############ DEBUG ############
test_input[32744:32751] = '{20.1317863606, 49.8565813904, 23.7659253278, -61.886236172, 42.8482103125, 6.17595155219, 2.85761979525, 33.323966411};
test_label[4093] = '{20.1317863606};
test_output[4093] = '{29.7256989676};
############ END DEBUG ############*/
test_input[32752:32759] = '{32'h4286ed91, 32'h42ac6e11, 32'h4265054a, 32'h414ccbf5, 32'hc2b76e0f, 32'hc113335d, 32'h42137678, 32'hc2365267};
test_label[4094] = '{32'h42137678};
test_output[4094] = '{32'h424565aa};
/*############ DEBUG ############
test_input[32752:32759] = '{67.4639970397, 86.2149727762, 57.2551656836, 12.7997942141, -91.7149566497, -9.20004013187, 36.8656931202, -45.5804710488};
test_label[4094] = '{36.8656931202};
test_output[4094] = '{49.3492796632};
############ END DEBUG ############*/
test_input[32760:32767] = '{32'hc2c56957, 32'h41f1b135, 32'hc211c37e, 32'hc204cb25, 32'hc2a03399, 32'hc0bd91cd, 32'hc1869fcf, 32'h419cd7d3};
test_label[4095] = '{32'hc211c37e};
test_output[4095] = '{32'h42854e10};
/*############ DEBUG ############
test_input[32760:32767] = '{-98.7057395775, 30.2115271316, -36.4409120444, -33.1983817312, -80.1007733967, -5.92404782557, -16.8280309105, 19.6053829231};
test_label[4095] = '{-36.4409120444};
test_output[4095] = '{66.6524639391};
############ END DEBUG ############*/
test_input[32768:32775] = '{32'h428e90c8, 32'h412981eb, 32'hc202a04c, 32'h4271bf13, 32'hc2b5d4ce, 32'hc0afe4b4, 32'hc2907ff5, 32'h42ac4db0};
test_label[4096] = '{32'hc202a04c};
test_output[4096] = '{32'h42ed9dd6};
/*############ DEBUG ############
test_input[32768:32775] = '{71.2827744752, 10.5942182493, -32.6565415494, 60.4365951523, -90.9156364547, -5.49666778704, -72.2499190231, 86.1517299018};
test_label[4096] = '{-32.6565415494};
test_output[4096] = '{118.8082718};
############ END DEBUG ############*/
test_input[32776:32783] = '{32'h42a6dde2, 32'h42189770, 32'h42b1226b, 32'hc13fcf11, 32'h4299171b, 32'h42ac4ca1, 32'hc1ed5011, 32'h42c78926};
test_label[4097] = '{32'h42c78926};
test_output[4097] = '{32'h377b0e14};
/*############ DEBUG ############
test_input[32776:32783] = '{83.43336699, 38.1478893849, 88.5672250896, -11.9880533049, 76.5451278563, 86.1496688476, -29.6640954623, 99.7678678599};
test_label[4097] = '{99.7678678599};
test_output[4097] = '{1.49640440581e-05};
############ END DEBUG ############*/
test_input[32784:32791] = '{32'h42016963, 32'hc2baa2a7, 32'h42b248a3, 32'hc244dd51, 32'h40a5306a, 32'h4282cc5c, 32'h4288bab2, 32'h4214d078};
test_label[4098] = '{32'h4282cc5c};
test_output[4098] = '{32'h41bdf11c};
/*############ DEBUG ############
test_input[32784:32791] = '{32.3529184186, -93.3176812953, 89.1418658946, -49.2161284692, 5.16215970204, 65.3991375767, 68.3646393513, 37.2035815834};
test_label[4098] = '{65.3991375767};
test_output[4098] = '{23.7427283189};
############ END DEBUG ############*/
test_input[32792:32799] = '{32'h429cac60, 32'h42c4a136, 32'h42b9a29a, 32'hc282f40b, 32'h424023a1, 32'h4155c097, 32'h42a234dc, 32'h42b1bb89};
test_label[4099] = '{32'h42b1bb89};
test_output[4099] = '{32'h41173e75};
/*############ DEBUG ############
test_input[32792:32799] = '{78.3366702287, 98.3148628806, 92.8175830875, -65.4766445684, 48.0347923361, 13.3595191774, 81.1032434272, 88.8662823097};
test_label[4099] = '{88.8662823097};
test_output[4099] = '{9.45274861292};
############ END DEBUG ############*/
test_input[32800:32807] = '{32'h42b31e7f, 32'h42612aec, 32'hc1c1a343, 32'hc288de9d, 32'hc2a52367, 32'hc2326dd2, 32'hc2bc4c92, 32'h423925c1};
test_label[4100] = '{32'h42b31e7f};
test_output[4100] = '{32'h27840000};
/*############ DEBUG ############
test_input[32800:32807] = '{89.5595594951, 56.2919171691, -24.2047176949, -68.4347927132, -82.5691431844, -44.6072465955, -94.1495482015, 46.2868676289};
test_label[4100] = '{89.5595594951};
test_output[4100] = '{3.66373598126e-15};
############ END DEBUG ############*/
test_input[32808:32815] = '{32'hc2858be4, 32'hc1b75973, 32'hc2c111be, 32'hc29d4466, 32'hc2b21886, 32'hc273706c, 32'h42979b0b, 32'hc21875a8};
test_label[4101] = '{32'hc2c111be};
test_output[4101] = '{32'h432c5664};
/*############ DEBUG ############
test_input[32808:32815] = '{-66.7732255709, -22.9186759337, -96.5346531653, -78.6335899057, -89.0478970607, -60.8597887715, 75.8028150722, -38.1148968905};
test_label[4101] = '{-96.5346531653};
test_output[4101] = '{172.337468238};
############ END DEBUG ############*/
test_input[32816:32823] = '{32'hc2b01e6d, 32'h42140fdf, 32'hc2b31b0a, 32'h4297fd4c, 32'hc219376c, 32'hc2a896db, 32'hc206ad9a, 32'hc1a76c75};
test_label[4102] = '{32'hc2b31b0a};
test_output[4102] = '{32'h43258c2b};
/*############ DEBUG ############
test_input[32816:32823] = '{-88.0594261341, 37.0154990736, -89.5528099503, 75.9947177968, -38.3041239582, -84.294642104, -33.6695344583, -20.92795842};
test_label[4102] = '{-89.5528099503};
test_output[4102] = '{165.547527747};
############ END DEBUG ############*/
test_input[32824:32831] = '{32'h42422b4e, 32'h418b703b, 32'hc2bf94ac, 32'hc22d8537, 32'h41ec7cb7, 32'h42b6e754, 32'hc2035e9d, 32'h4210fe02};
test_label[4103] = '{32'h42422b4e};
test_output[4103] = '{32'h422ba35a};
/*############ DEBUG ############
test_input[32824:32831] = '{48.5422902255, 17.4298000944, -95.7903752158, -43.3800930133, 29.56089603, 91.4518129515, -32.8423969802, 36.248054523};
test_label[4103] = '{48.5422902255};
test_output[4103] = '{42.909522726};
############ END DEBUG ############*/
test_input[32832:32839] = '{32'h4241dfff, 32'h411756c0, 32'hc26bf63b, 32'hc2bc5070, 32'hc18c0ad8, 32'h42457d7a, 32'hc2ac7ba8, 32'hc2baa332};
test_label[4104] = '{32'h4241dfff};
test_output[4104] = '{32'h3f9f3663};
/*############ DEBUG ############
test_input[32832:32839] = '{48.4687475324, 9.45867908326, -58.9904607307, -94.1571013393, -17.5052946395, 49.3725339207, -86.2415148778, -93.3187387702};
test_label[4104] = '{48.4687475324};
test_output[4104] = '{1.24384727791};
############ END DEBUG ############*/
test_input[32840:32847] = '{32'hc177707c, 32'h41ed9dca, 32'hc1d6d327, 32'hc21a0987, 32'h4235eccb, 32'hc2a27254, 32'hc2bd9804, 32'h42783168};
test_label[4105] = '{32'hc2a27254};
test_output[4105] = '{32'h430f4584};
/*############ DEBUG ############
test_input[32840:32847] = '{-15.464961599, 29.7020458232, -26.8531013136, -38.5093057743, 45.481243851, -81.2232981974, -94.7969052071, 62.0482496988};
test_label[4105] = '{-81.2232981974};
test_output[4105] = '{143.27154796};
############ END DEBUG ############*/
test_input[32848:32855] = '{32'h424bb46a, 32'hc2980646, 32'h42b1547f, 32'hc1017368, 32'h423b284c, 32'h41ad1f96, 32'h40f36827, 32'hc1dd58e1};
test_label[4106] = '{32'h42b1547f};
test_output[4106] = '{32'h80000000};
/*############ DEBUG ############
test_input[32848:32855] = '{50.9261860754, -76.0122505866, 88.6650336819, -8.09067516546, 46.7893514317, 21.6404219565, 7.60646396416, -27.6683973133};
test_label[4106] = '{88.6650336819};
test_output[4106] = '{-0.0};
############ END DEBUG ############*/
test_input[32856:32863] = '{32'h41b39753, 32'h4260ddd0, 32'hc2a7e391, 32'hc2143fc9, 32'hc2b28e7f, 32'hc275aa89, 32'h425f0bd0, 32'hc1c9a928};
test_label[4107] = '{32'hc2a7e391};
test_output[4107] = '{32'h430ca701};
/*############ DEBUG ############
test_input[32856:32863] = '{22.4488885071, 56.2166151237, -83.9444633138, -37.0622892608, -89.2783146404, -61.4165400308, 55.7615364151, -25.2075954998};
test_label[4107] = '{-83.9444633138};
test_output[4107] = '{140.652352999};
############ END DEBUG ############*/
test_input[32864:32871] = '{32'hc2a129a9, 32'hc207b485, 32'hc2326e3a, 32'h4271fb87, 32'hc27c5af2, 32'h42bdf834, 32'h419b9452, 32'hc22b0637};
test_label[4108] = '{32'hc2a129a9};
test_output[4108] = '{32'h432f90ee};
/*############ DEBUG ############
test_input[32864:32871] = '{-80.5813655889, -33.9262871856, -44.6076415608, 60.4956313156, -63.0888146355, 94.9847722919, 19.4474226487, -42.7560709438};
test_label[4108] = '{-80.5813655889};
test_output[4108] = '{175.566137881};
############ END DEBUG ############*/
test_input[32872:32879] = '{32'h4171c255, 32'h428195e6, 32'h42982fbf, 32'hc22ae509, 32'h427c572f, 32'hc2307b57, 32'hc095f04f, 32'hc227372b};
test_label[4109] = '{32'hc227372b};
test_output[4109] = '{32'h42ebcb56};
/*############ DEBUG ############
test_input[32872:32879] = '{15.1099447555, 64.7927741632, 76.0932526214, -42.7236658037, 63.0851405421, -44.1204472446, -4.68558441724, -41.8038757369};
test_label[4109] = '{-41.8038757369};
test_output[4109] = '{117.897142967};
############ END DEBUG ############*/
test_input[32880:32887] = '{32'h41991207, 32'hc2b478f7, 32'h4268b799, 32'hc2781907, 32'h4122d51c, 32'h414dcd62, 32'hbf35a36f, 32'hc2897948};
test_label[4110] = '{32'h414dcd62};
test_output[4110] = '{32'h42354441};
/*############ DEBUG ############
test_input[32880:32887] = '{19.1338032253, -90.2362559684, 58.1792954382, -62.0244425428, 10.177028787, 12.8626427345, -0.709525036245, -68.7368806124};
test_label[4110] = '{12.8626427345};
test_output[4110] = '{45.3166527037};
############ END DEBUG ############*/
test_input[32888:32895] = '{32'h42aebb1b, 32'h429581d7, 32'h4246f895, 32'hc23a736f, 32'h42786db2, 32'h41d472f7, 32'h4253252c, 32'hc243b126};
test_label[4111] = '{32'h429581d7};
test_output[4111] = '{32'h4149ca2a};
/*############ DEBUG ############
test_input[32888:32895] = '{87.3654440395, 74.7535913072, 49.7427571714, -46.6127285728, 62.1071258935, 26.5561344235, 52.7863017726, -48.9229951663};
test_label[4111] = '{74.7535913072};
test_output[4111] = '{12.6118560646};
############ END DEBUG ############*/
test_input[32896:32903] = '{32'hc24a2017, 32'hc27a818e, 32'h42824830, 32'h42a167cf, 32'hc2506a34, 32'hc2c5fbc4, 32'h42ba90c3, 32'h4155ad46};
test_label[4112] = '{32'h42ba90c3};
test_output[4112] = '{32'h3666dded};
/*############ DEBUG ############
test_input[32896:32903] = '{-50.5313372103, -62.626516628, 65.1409932977, 80.7027546523, -52.103715317, -98.9917281037, 93.2827384627, 13.354802973};
test_label[4112] = '{93.2827384627};
test_output[4112] = '{3.44018483794e-06};
############ END DEBUG ############*/
test_input[32904:32911] = '{32'hc2b1e254, 32'hc2b458e2, 32'hc2854b11, 32'h40f496c8, 32'hc2625114, 32'h409890da, 32'hc2b8958e, 32'h3f6551e9};
test_label[4113] = '{32'hc2854b11};
test_output[4113] = '{32'h4294b123};
/*############ DEBUG ############
test_input[32904:32911] = '{-88.9420503935, -90.1735998037, -66.6466108195, 7.64340588165, -56.5791779767, 4.7676821535, -92.292097799, 0.89578108646};
test_label[4113] = '{-66.6466108195};
test_output[4113] = '{74.3459706566};
############ END DEBUG ############*/
test_input[32912:32919] = '{32'h42959da7, 32'hc28eb4ad, 32'h421f77fd, 32'h4253c0ee, 32'h4257c1ba, 32'h41814ad3, 32'hc0edc5e2, 32'h42afca63};
test_label[4114] = '{32'h4253c0ee};
test_output[4114] = '{32'h420bd3d9};
/*############ DEBUG ############
test_input[32912:32919] = '{74.8079116294, -71.3528847318, 39.8671761227, 52.9384067055, 53.9391860002, 16.1615358393, -7.43040568052, 87.8952873531};
test_label[4114] = '{52.9384067055};
test_output[4114] = '{34.9568827189};
############ END DEBUG ############*/
test_input[32920:32927] = '{32'h4256cf64, 32'h4281520e, 32'hc2a47c6e, 32'h429d8a13, 32'h42349ba1, 32'hc2be3274, 32'hc200bee1, 32'h42ba8139};
test_label[4115] = '{32'h429d8a13};
test_output[4115] = '{32'h4167b932};
/*############ DEBUG ############
test_input[32920:32927] = '{53.7025317342, 64.6602618464, -82.2430293099, 78.7696727785, 45.1519831131, -95.098538356, -32.1864037675, 93.2523855044};
test_label[4115] = '{78.7696727785};
test_output[4115] = '{14.4827132391};
############ END DEBUG ############*/
test_input[32928:32935] = '{32'hc2802a6e, 32'hc2a107f6, 32'hc1eca952, 32'h4281d2fa, 32'h4093a7fd, 32'hc2a99701, 32'h42b779e8, 32'hc0d0e194};
test_label[4116] = '{32'hc2802a6e};
test_output[4116] = '{32'h431bd22b};
/*############ DEBUG ############
test_input[32928:32935] = '{-64.0828668948, -80.5155476395, -29.5826765064, 64.9120657606, 4.61425631788, -84.7949294974, 91.7380984243, -6.52753623144};
test_label[4116] = '{-64.0828668948};
test_output[4116] = '{155.820965319};
############ END DEBUG ############*/
test_input[32936:32943] = '{32'hc2315169, 32'hc14f205b, 32'h4259a4c8, 32'h428e858b, 32'hc226c1dc, 32'hc291f47c, 32'h40ecc876, 32'hc1f801ef};
test_label[4117] = '{32'hc226c1dc};
test_output[4117] = '{32'h42e1e67a};
/*############ DEBUG ############
test_input[32936:32943] = '{-44.3295034447, -12.9453992627, 54.4109209069, 71.2608290247, -41.6893170106, -72.9775114577, 7.39947016446, -31.0009447856};
test_label[4117] = '{-41.6893170106};
test_output[4117] = '{112.950146083};
############ END DEBUG ############*/
test_input[32944:32951] = '{32'hc097d6bd, 32'h42813ac7, 32'h42797240, 32'hc2c2eba3, 32'h422d019e, 32'hc28a232e, 32'hc2bc7d17, 32'h42a5bf31};
test_label[4118] = '{32'hc2c2eba3};
test_output[4118] = '{32'h4334556a};
/*############ DEBUG ############
test_input[32944:32951] = '{-4.74496293806, 64.6148028387, 62.3615705114, -97.4602253335, 43.2515784856, -69.0687121396, -94.244312396, 82.8734186436};
test_label[4118] = '{-97.4602253335};
test_output[4118] = '{180.33364399};
############ END DEBUG ############*/
test_input[32952:32959] = '{32'h42bb882e, 32'hc2795bd1, 32'h40afea5b, 32'h42031506, 32'hc1dd060e, 32'h42b88efc, 32'hc20df6bb, 32'h41c162bd};
test_label[4119] = '{32'h41c162bd};
test_output[4119] = '{32'h428b97de};
/*############ DEBUG ############
test_input[32952:32959] = '{93.7659770568, -62.3396626959, 5.4973578174, 32.7705296617, -27.6279564654, 92.2792700845, -35.4909476203, 24.1732119852};
test_label[4119] = '{24.1732119852};
test_output[4119] = '{69.7966165517};
############ END DEBUG ############*/
test_input[32960:32967] = '{32'h42ab8228, 32'hc19d4083, 32'hc243355f, 32'h421cc4cc, 32'hc113d893, 32'hc26cdf3b, 32'h412909f1, 32'h425bac14};
test_label[4120] = '{32'hc19d4083};
test_output[4120] = '{32'h42d2d249};
/*############ DEBUG ############
test_input[32960:32967] = '{85.7542148972, -19.6565000548, -48.8021210008, 39.1921842408, -9.24037478418, -59.2179993726, 10.5649271075, 54.9180449351};
test_label[4120] = '{-19.6565000548};
test_output[4120] = '{105.410714952};
############ END DEBUG ############*/
test_input[32968:32975] = '{32'hc2925d44, 32'hc1964287, 32'h42333ee2, 32'hc2b9662a, 32'h42194977, 32'h4246bc25, 32'h40a1dda7, 32'hc18f8591};
test_label[4121] = '{32'hc2b9662a};
test_output[4121] = '{32'h430e6412};
/*############ DEBUG ############
test_input[32968:32975] = '{-73.1821632147, -18.782484729, 44.8114078323, -92.6995361812, 38.3217445216, 49.6837330291, 5.05830730767, -17.9402176239};
test_label[4121] = '{-92.6995361812};
test_output[4121] = '{142.39090714};
############ END DEBUG ############*/
test_input[32976:32983] = '{32'hc185cf1c, 32'h42116b49, 32'h42b2d7ed, 32'h42a1ff63, 32'h42b3e89b, 32'h42b5426b, 32'h428cf170, 32'h41f018a1};
test_label[4122] = '{32'h42b3e89b};
test_output[4122] = '{32'h3fa23e66};
/*############ DEBUG ############
test_input[32976:32983] = '{-16.7261274304, 36.3547707813, 89.4217299209, 80.9987993947, 89.9543104645, 90.6297254878, 70.4715594747, 30.0120255766};
test_label[4122] = '{89.9543104645};
test_output[4122] = '{1.26752920875};
############ END DEBUG ############*/
test_input[32984:32991] = '{32'h4207cb2a, 32'hc2b05c95, 32'h429897f4, 32'h420dc1ce, 32'h420c7a62, 32'hc220733d, 32'hc2ba0499, 32'hc248c28b};
test_label[4123] = '{32'h420c7a62};
test_output[4123] = '{32'h4224b586};
/*############ DEBUG ############
test_input[32984:32991] = '{33.948402774, -88.1808228011, 76.2967824124, 35.439262999, 35.1195133024, -40.1125362011, -93.0089782803, -50.1899831517};
test_label[4123] = '{35.1195133024};
test_output[4123] = '{41.17726911};
############ END DEBUG ############*/
test_input[32992:32999] = '{32'hc22223e8, 32'hc1cb35a8, 32'h419ee7f5, 32'h429d2048, 32'h41863561, 32'hc2c06a09, 32'h4290b894, 32'h42986efe};
test_label[4124] = '{32'hc1cb35a8};
test_output[4124] = '{32'h42d01d72};
/*############ DEBUG ############
test_input[32992:32999] = '{-40.5350662044, -25.401199421, 19.8632606215, 78.5630455405, 16.7760642358, -96.2071023368, 72.3605046944, 76.2167807908};
test_label[4124] = '{-25.401199421};
test_output[4124] = '{104.057507899};
############ END DEBUG ############*/
test_input[33000:33007] = '{32'h40953b7e, 32'h40ce4e26, 32'h42a4523b, 32'hc1e740a4, 32'h40af9b63, 32'h4215e553, 32'hc1d2d880, 32'h422eb3de};
test_label[4125] = '{32'hc1d2d880};
test_output[4125] = '{32'h42d9085b};
/*############ DEBUG ############
test_input[33000:33007] = '{4.6635123241, 6.44703969704, 82.1606095252, -28.9065633827, 5.48771814188, 37.4739491581, -26.3557131452, 43.6756502076};
test_label[4125] = '{-26.3557131452};
test_output[4125] = '{108.51632267};
############ END DEBUG ############*/
test_input[33008:33015] = '{32'h425c87db, 32'hc2a0835a, 32'hc25feb4a, 32'h4256e542, 32'hc2706cc9, 32'hc2639025, 32'hc2a9df55, 32'h40824357};
test_label[4126] = '{32'hc2706cc9};
test_output[4126] = '{32'h42e6ea4a};
/*############ DEBUG ############
test_input[33008:33015] = '{55.1326715119, -80.2565490654, -55.9797759184, 53.7238853016, -60.106237233, -56.8907670408, -84.9361937591, 4.07071998752};
test_label[4126] = '{-60.106237233};
test_output[4126] = '{115.457594215};
############ END DEBUG ############*/
test_input[33016:33023] = '{32'hc274a50a, 32'hc1091bda, 32'hc1b4f8b0, 32'h42b8cc8e, 32'h41a32d80, 32'h424a5d39, 32'h4226d6af, 32'h420e959a};
test_label[4127] = '{32'hc1b4f8b0};
test_output[4127] = '{32'h42e60aba};
/*############ DEBUG ############
test_input[33016:33023] = '{-61.1611721569, -8.56929951712, -22.6214296738, 92.3995194094, 20.3972159677, 50.5910375066, 41.7096514655, 35.6460934633};
test_label[4127] = '{-22.6214296738};
test_output[4127] = '{115.020949083};
############ END DEBUG ############*/
test_input[33024:33031] = '{32'h42a46541, 32'hc2b501c6, 32'h422fa2b9, 32'hc25dc6df, 32'h3fa40f87, 32'h40119fdd, 32'h4268c985, 32'hc2b3259b};
test_label[4128] = '{32'hc2b501c6};
test_output[4128] = '{32'h432cb384};
/*############ DEBUG ############
test_input[33024:33031] = '{82.1977620088, -90.5034643668, 43.9089074529, -55.444208643, 1.28172383027, 2.27538225554, 58.1967955987, -89.5734503088};
test_label[4128] = '{-90.5034643668};
test_output[4128] = '{172.701226376};
############ END DEBUG ############*/
test_input[33032:33039] = '{32'h4295446a, 32'h42aec528, 32'hc284deed, 32'h41e43676, 32'hc1faa0a7, 32'h424e5b3f, 32'hbf89c0e2, 32'h40e5379a};
test_label[4129] = '{32'h4295446a};
test_output[4129] = '{32'h414c05ef};
/*############ DEBUG ############
test_input[33032:33039] = '{74.6336237667, 87.385069874, -66.435405435, 28.5265918968, -31.3284433902, 51.5891063634, -1.07619880856, 7.16303725068};
test_label[4129] = '{74.6336237667};
test_output[4129] = '{12.7514490055};
############ END DEBUG ############*/
test_input[33040:33047] = '{32'h41bf63bd, 32'h4274b07f, 32'h4134c6e5, 32'hc1a25b62, 32'hc2583044, 32'h42b40d0b, 32'h3f527198, 32'hc25a7f99};
test_label[4130] = '{32'h4134c6e5};
test_output[4130] = '{32'h429d742e};
/*############ DEBUG ############
test_input[33040:33047] = '{23.923700083, 61.1723603735, 11.2985584956, -20.294620397, -54.0471326096, 90.0254743173, 0.822045776355, -54.6246051886};
test_label[4130] = '{11.2985584956};
test_output[4130] = '{78.7269158217};
############ END DEBUG ############*/
test_input[33048:33055] = '{32'h41cb460a, 32'h429b481b, 32'hc23873af, 32'h41aa5f73, 32'h4276e220, 32'h42587a31, 32'h428f9cb1, 32'h40b88929};
test_label[4131] = '{32'h42587a31};
test_output[4131] = '{32'h41bc3205};
/*############ DEBUG ############
test_input[33048:33055] = '{25.4091996104, 77.6408308785, -46.1129707428, 21.2966064439, 61.7208234644, 54.1193262644, 71.8060379668, 5.76674321118};
test_label[4131] = '{54.1193262644};
test_output[4131] = '{23.5244244977};
############ END DEBUG ############*/
test_input[33056:33063] = '{32'h429c5144, 32'hc235dcf5, 32'hc287ff4c, 32'h417380e3, 32'hc24f79fd, 32'hc2447b14, 32'h42a5f122, 32'hc29a5933};
test_label[4132] = '{32'hc29a5933};
test_output[4132] = '{32'h4320273d};
/*############ DEBUG ############
test_input[33056:33063] = '{78.1587244703, -45.4657798985, -67.9986305192, 15.2189668529, -51.8691289535, -49.1201923522, 82.9709617196, -77.1742154652};
test_label[4132] = '{-77.1742154652};
test_output[4132] = '{160.153273968};
############ END DEBUG ############*/
test_input[33064:33071] = '{32'hc2596f4b, 32'hc23dcb04, 32'h4261a8c5, 32'h41a4b8d6, 32'h41603cbe, 32'h42b5415d, 32'hc10dce67, 32'h42aa966c};
test_label[4133] = '{32'h42b5415d};
test_output[4133] = '{32'h3b9dbcaf};
/*############ DEBUG ############
test_input[33064:33071] = '{-54.3586832541, -47.4482583324, 56.4148149913, 20.5902516054, 14.0148300616, 90.6276645014, -8.86289132385, 85.2937940345};
test_label[4133] = '{90.6276645014};
test_output[4133] = '{0.00481375271519};
############ END DEBUG ############*/
test_input[33072:33079] = '{32'hc1a06359, 32'h42b71175, 32'hc271bff2, 32'hc23859fa, 32'h41a86561, 32'h42a26ebd, 32'h42b1084f, 32'h42a49a26};
test_label[4134] = '{32'hc23859fa};
test_output[4134] = '{32'h4309ab7a};
/*############ DEBUG ############
test_input[33072:33079] = '{-20.0485095598, 91.5340960948, -60.4374451753, -46.0878665092, 21.0495010085, 81.2162858469, 88.5162278063, 82.3010701951};
test_label[4134] = '{-46.0878665092};
test_output[4134] = '{137.6698344};
############ END DEBUG ############*/
test_input[33080:33087] = '{32'h4200ad30, 32'h42514e1e, 32'h42b7ea09, 32'h42b9d3eb, 32'hc265d167, 32'hc2b93774, 32'hc214389f, 32'h41be175c};
test_label[4135] = '{32'hc214389f};
test_output[4135] = '{32'h43024b55};
/*############ DEBUG ############
test_input[33080:33087] = '{32.1691299446, 52.3262857048, 91.9571035819, 92.9138995659, -57.4544948353, -92.6083080116, -37.0552953985, 23.7614068302};
test_label[4135] = '{-37.0552953985};
test_output[4135] = '{130.294260714};
############ END DEBUG ############*/
test_input[33088:33095] = '{32'hc204af5f, 32'hc28c3444, 32'hc294bc7b, 32'h42483e5d, 32'h4241d051, 32'h40ff9090, 32'h424efc71, 32'h42c238c2};
test_label[4136] = '{32'h42c238c2};
test_output[4136] = '{32'h80000000};
/*############ DEBUG ############
test_input[33088:33095] = '{-33.1712600368, -70.102081934, -74.3681259844, 50.0609016694, 48.4534357684, 7.98639657347, 51.7465247162, 97.1108541782};
test_label[4136] = '{97.1108541782};
test_output[4136] = '{-0.0};
############ END DEBUG ############*/
test_input[33096:33103] = '{32'h424537e0, 32'h429909ce, 32'h42aed8ba, 32'h42b6ea9b, 32'h42543cd6, 32'hc2b1729b, 32'hc1e236e1, 32'hc2b4dd38};
test_label[4137] = '{32'hc1e236e1};
test_output[4137] = '{32'h42ef814d};
/*############ DEBUG ############
test_input[33096:33103] = '{49.3045669969, 76.5191508651, 87.4232976327, 91.4582148328, 53.0594117957, -88.7238412799, -28.2767962288, -90.4320655715};
test_label[4137] = '{-28.2767962288};
test_output[4137] = '{119.752543928};
############ END DEBUG ############*/
test_input[33104:33111] = '{32'h4154fa67, 32'h4201c7a9, 32'h42bae1e7, 32'hc2816ca2, 32'h423e981b, 32'hc21272fb, 32'hc29d437e, 32'hc29e5786};
test_label[4138] = '{32'h4201c7a9};
test_output[4138] = '{32'h4273fc25};
/*############ DEBUG ############
test_input[33104:33111] = '{13.3111330505, 32.4449788107, 93.4412155603, -64.7121716975, 47.6485417629, -36.612284076, -78.6318181896, -79.1709458647};
test_label[4138] = '{32.4449788107};
test_output[4138] = '{60.9962367496};
############ END DEBUG ############*/
test_input[33112:33119] = '{32'h413f5839, 32'h42ad7b7f, 32'h417b0a66, 32'h40160378, 32'hc29790e5, 32'h416190cf, 32'hc1bd0ea6, 32'hc28e377f};
test_label[4139] = '{32'h413f5839};
test_output[4139] = '{32'h42959078};
/*############ DEBUG ############
test_input[33112:33119] = '{11.9590382638, 86.7412055813, 15.6900389376, 2.34396173071, -75.7829998693, 14.0978536934, -23.632153233, -71.1083937046};
test_label[4139] = '{11.9590382638};
test_output[4139] = '{74.7821673175};
############ END DEBUG ############*/
test_input[33120:33127] = '{32'hbfcc567d, 32'h42a33cf3, 32'hc21b64ae, 32'hc28696ea, 32'hc25fb4f9, 32'h42b8a208, 32'h40f3541f, 32'hc0b6933a};
test_label[4140] = '{32'h40f3541f};
test_output[4140] = '{32'h42a96cc9};
/*############ DEBUG ############
test_input[33120:33127] = '{-1.59638943001, 81.6190420259, -38.8483202683, -67.2947532881, -55.9267304334, 92.3164691198, 7.60401846642, -5.70547195345};
test_label[4140] = '{7.60401846642};
test_output[4140] = '{84.7124732561};
############ END DEBUG ############*/
test_input[33128:33135] = '{32'hc29d32c9, 32'hc2c1fa00, 32'h428d0b34, 32'hc28f8466, 32'hc2c7d211, 32'h42a0af06, 32'hc265a49c, 32'hc2189a96};
test_label[4141] = '{32'hc2c1fa00};
test_output[4141] = '{32'h43315487};
/*############ DEBUG ############
test_input[33128:33135] = '{-78.5991881974, -96.9882812488, 70.5218790618, -71.7585881153, -99.9102879566, 80.3418441265, -57.4107511709, -38.150961995};
test_label[4141] = '{-96.9882812488};
test_output[4141] = '{177.330179729};
############ END DEBUG ############*/
test_input[33136:33143] = '{32'hc2c58aba, 32'hc15419d5, 32'hc2666299, 32'h42873ebc, 32'h42c4dce0, 32'hc1dded6e, 32'hc1ce9cb6, 32'hc299da0e};
test_label[4142] = '{32'hc15419d5};
test_output[4142] = '{32'h42df601b};
/*############ DEBUG ############
test_input[33136:33143] = '{-98.7709500957, -13.256306772, -57.5962855459, 67.6225295599, 98.4313956159, -27.7409328455, -25.8265195009, -76.9258871186};
test_label[4142] = '{-13.256306772};
test_output[4142] = '{111.687702388};
############ END DEBUG ############*/
test_input[33144:33151] = '{32'hc1eca142, 32'h429cfd55, 32'h42bbddd7, 32'h42b1cfd5, 32'h421277ec, 32'h42332db7, 32'hc297fc13, 32'hc29e8390};
test_label[4143] = '{32'h42b1cfd5};
test_output[4143] = '{32'h40a115b6};
/*############ DEBUG ############
test_input[33144:33151] = '{-29.5787383106, 78.4947895363, 93.9332836447, 88.9059184764, 36.6171118748, 44.7946422456, -75.992332191, -79.2569571426};
test_label[4143] = '{88.9059184764};
test_output[4143] = '{5.03390002874};
############ END DEBUG ############*/
test_input[33152:33159] = '{32'h427d5cdf, 32'hc1909905, 32'h428e68a4, 32'hc280d439, 32'hc19d1f16, 32'h418c2876, 32'hc24be3f1, 32'hc11b32a4};
test_label[4144] = '{32'hc280d439};
test_output[4144] = '{32'h43079e88};
/*############ DEBUG ############
test_input[33152:33159] = '{63.340695654, -18.074717245, 71.2043777058, -64.4144947897, -19.6401788348, 17.5197565078, -50.972598884, -9.69986371697};
test_label[4144] = '{-64.4144947897};
test_output[4144] = '{135.619256877};
############ END DEBUG ############*/
test_input[33160:33167] = '{32'hc2430fda, 32'h42a0e021, 32'h429b60e7, 32'hc22c64a7, 32'h4204a460, 32'h4255e8c1, 32'h40f4f9a2, 32'h428cb71c};
test_label[4145] = '{32'h42a0e021};
test_output[4145] = '{32'h3d7e5a35};
/*############ DEBUG ############
test_input[33160:33167] = '{-48.7654818836, 80.4377527906, 77.6892624479, -43.0982924569, 33.160522674, 53.4772969674, 7.65547274256, 70.3576370194};
test_label[4145] = '{80.4377527906};
test_output[4145] = '{0.0620977459505};
############ END DEBUG ############*/
test_input[33168:33175] = '{32'h419ac62a, 32'h428153c7, 32'h425dceda, 32'h4270fa6f, 32'h3fb41df3, 32'h4238dc24, 32'hc2863838, 32'h4276466f};
test_label[4146] = '{32'hc2863838};
test_output[4146] = '{32'h4303d44b};
/*############ DEBUG ############
test_input[33168:33175] = '{19.3467598008, 64.6636258942, 55.4520018616, 60.2445621644, 1.40716395029, 46.2149806776, -67.1098029063, 61.5687824422};
test_label[4146] = '{-67.1098029063};
test_output[4146] = '{131.82926786};
############ END DEBUG ############*/
test_input[33176:33183] = '{32'h4257db41, 32'hc256a85d, 32'hc20260c3, 32'h40f1fdc4, 32'h41e175a6, 32'h42b5e608, 32'h42b5fbfc, 32'hc2897a12};
test_label[4147] = '{32'h4257db41};
test_output[4147] = '{32'h4216ccc8};
/*############ DEBUG ############
test_input[33176:33183] = '{53.9641137108, -53.6644176645, -32.5944930636, 7.56222740314, 28.1824451176, 90.9492809775, 90.9921544083, -68.7384195231};
test_label[4147] = '{53.9641137108};
test_output[4147] = '{37.6999809114};
############ END DEBUG ############*/
test_input[33184:33191] = '{32'h42bf67d5, 32'h420d1d1a, 32'hc1afdf9b, 32'h42a0c5a6, 32'hc27a7193, 32'hc2a1f45f, 32'hc2bc4fdf, 32'h42bc3e80};
test_label[4148] = '{32'h42a0c5a6};
test_output[4148] = '{32'h41781019};
/*############ DEBUG ############
test_input[33184:33191] = '{95.7027990633, 35.2784205912, -21.9841832967, 80.38603372, -62.6109114083, -80.9772883005, -94.1559949638, 94.1220740352};
test_label[4148] = '{80.38603372};
test_output[4148] = '{15.5039301836};
############ END DEBUG ############*/
test_input[33192:33199] = '{32'hc27e9c6b, 32'hc1905ba8, 32'hc103bf16, 32'h40804e4d, 32'h42ab9fcf, 32'hc23c8aca, 32'h41706bee, 32'hc1ad9273};
test_label[4149] = '{32'h40804e4d};
test_output[4149] = '{32'h42a39aea};
/*############ DEBUG ############
test_input[33192:33199] = '{-63.6527508765, -18.0447546869, -8.23415204717, 4.00955838716, 85.8121234615, -47.1355347853, 15.0263504288, -21.6965082751};
test_label[4149] = '{4.00955838716};
test_output[4149] = '{81.8025650744};
############ END DEBUG ############*/
test_input[33200:33207] = '{32'h424cb276, 32'h41b138ce, 32'hc1f8a75e, 32'h41f52cfd, 32'h42aee1ea, 32'hc2039379, 32'h42c75475, 32'h42bb7160};
test_label[4150] = '{32'h42c75475};
test_output[4150] = '{32'h3b2bfb5c};
/*############ DEBUG ############
test_input[33200:33207] = '{51.1742800032, 22.1527367231, -31.0817213095, 30.6469666148, 87.4412382543, -32.8940166764, 99.664958258, 93.7214335341};
test_label[4150] = '{99.664958258};
test_output[4150] = '{0.00262423502214};
############ END DEBUG ############*/
test_input[33208:33215] = '{32'h429bbacc, 32'h40d2f092, 32'hc2073132, 32'hc27818f6, 32'hc23de7e8, 32'hc23a5667, 32'h423d053a, 32'h41ece93f};
test_label[4151] = '{32'hc23a5667};
test_output[4151] = '{32'h42f8e600};
/*############ DEBUG ############
test_input[33208:33215] = '{77.8648381682, 6.59186641625, -33.7980410188, -62.02437742, -47.4764713782, -46.5843784137, 47.2551021703, 29.6138890051};
test_label[4151] = '{-46.5843784137};
test_output[4151] = '{124.449216582};
############ END DEBUG ############*/
test_input[33216:33223] = '{32'hc0ffb708, 32'h41cbe1db, 32'hc1293ebc, 32'h42a3f1ac, 32'h4108e010, 32'h417fe412, 32'hc1b77966, 32'h4222989a};
test_label[4152] = '{32'hc1293ebc};
test_output[4152] = '{32'h42b91984};
/*############ DEBUG ############
test_input[33216:33223] = '{-7.99109261139, 25.4852811107, -10.5778157575, 81.97201639, 8.55470273595, 15.9931813567, -22.9342774105, 40.6490252852};
test_label[4152] = '{-10.5778157575};
test_output[4152] = '{92.5498321475};
############ END DEBUG ############*/
test_input[33224:33231] = '{32'hc231d6d7, 32'hc2c5801a, 32'h428d0f10, 32'h420c7e8e, 32'h42c0030b, 32'hbfcb4a6a, 32'h420ba2fb, 32'hc2c59e6d};
test_label[4153] = '{32'h428d0f10};
test_output[4153] = '{32'h41cbcfe9};
/*############ DEBUG ############
test_input[33224:33231] = '{-44.4598056827, -98.7501948145, 70.5294216923, 35.1235883793, 96.0059394855, -1.5882084898, 34.909159771, -98.809425886};
test_label[4153] = '{70.5294216923};
test_output[4153] = '{25.4765177932};
############ END DEBUG ############*/
test_input[33232:33239] = '{32'hc0f53744, 32'hc006af06, 32'h41478523, 32'h4283017a, 32'h42b18565, 32'hc1e06eac, 32'hc2a8fe7b, 32'hc29d6ec7};
test_label[4154] = '{32'h41478523};
test_output[4154] = '{32'h429894c1};
/*############ DEBUG ############
test_input[33232:33239] = '{-7.66299623953, -2.10443261741, 12.4700042916, 65.5028836714, 88.7605364766, -28.0540398327, -84.4970352148, -78.7163615492};
test_label[4154] = '{12.4700042916};
test_output[4154] = '{76.2905321851};
############ END DEBUG ############*/
test_input[33240:33247] = '{32'hc29f4065, 32'h42b281f3, 32'hc2abcc8b, 32'hc288400e, 32'h42908df3, 32'h3fe5b47d, 32'hc27121bd, 32'hc2914523};
test_label[4155] = '{32'hc27121bd};
test_output[4155] = '{32'h43158969};
/*############ DEBUG ############
test_input[33240:33247] = '{-79.6257683995, 89.2538077377, -85.899498551, -68.1251043093, 72.2772450527, 1.79457052225, -60.282948235, -72.6350344103};
test_label[4155] = '{-60.282948235};
test_output[4155] = '{149.536756015};
############ END DEBUG ############*/
test_input[33248:33255] = '{32'hc2c32803, 32'h419e189e, 32'hc1084115, 32'hbfffc8e9, 32'hc2544bd6, 32'hc14af655, 32'hc20b7515, 32'hc271442f};
test_label[4156] = '{32'hc2544bd6};
test_output[4156] = '{32'h4291ac12};
/*############ DEBUG ############
test_input[33248:33255] = '{-97.5781453437, 19.7620202767, -8.51588945684, -1.99831875796, -53.0740574276, -12.6851392222, -34.8643381705, -60.3165845568};
test_label[4156] = '{-53.0740574276};
test_output[4156] = '{72.8360777047};
############ END DEBUG ############*/
test_input[33256:33263] = '{32'h4256c25a, 32'hc29240c7, 32'h4117b0d0, 32'hc1f0d116, 32'h4191fcc8, 32'hc2a04676, 32'hc1d8bd06, 32'hc20cea00};
test_label[4157] = '{32'hc20cea00};
test_output[4157] = '{32'h42b1d62d};
/*############ DEBUG ############
test_input[33256:33263] = '{53.6897947997, -73.1265215448, 9.48066745224, -30.1020921665, 18.2484289597, -80.1376182914, -27.0922975227, -35.2285153092};
test_label[4157] = '{-35.2285153092};
test_output[4157] = '{88.9183101089};
############ END DEBUG ############*/
test_input[33264:33271] = '{32'h41621a29, 32'hc2a1df4a, 32'hc148adca, 32'h41f44e11, 32'hc28f23ad, 32'h42392485, 32'hc2320e29, 32'hc195df75};
test_label[4158] = '{32'h41621a29};
test_output[4158] = '{32'h42009dfb};
/*############ DEBUG ############
test_input[33264:33271] = '{14.1313864587, -80.9361102948, -12.5424286839, 30.5381184607, -71.5696826057, 46.2856643315, -44.5138275269, -18.7341107133};
test_label[4158] = '{14.1313864587};
test_output[4158] = '{32.1542780176};
############ END DEBUG ############*/
test_input[33272:33279] = '{32'hc2ba35c1, 32'hc1a01f7f, 32'h42a3b84d, 32'hc2b65d3c, 32'hc19dc95c, 32'hc1c40f30, 32'h41579071, 32'hc2c1baf5};
test_label[4159] = '{32'h41579071};
test_output[4159] = '{32'h4288c63f};
/*############ DEBUG ############
test_input[33272:33279] = '{-93.1049867003, -20.015378636, 81.8599625812, -91.1820966778, -19.7233192957, -24.5074166484, 13.4727640168, -96.865151211};
test_label[4159] = '{13.4727640168};
test_output[4159] = '{68.3871985644};
############ END DEBUG ############*/
test_input[33280:33287] = '{32'hc2164280, 32'h41f3d2ef, 32'h4263da4b, 32'hc18aad7c, 32'h429012f5, 32'h40c375c3, 32'h420213ea, 32'hc286af6a};
test_label[4160] = '{32'h4263da4b};
test_output[4160] = '{32'h41712e7f};
/*############ DEBUG ############
test_input[33280:33287] = '{-37.5649399035, 30.4779949208, 56.9631777761, -17.3347099544, 72.037028734, 6.10812511145, 32.5194481635, -67.3426086781};
test_label[4160] = '{56.9631777761};
test_output[4160] = '{15.073851242};
############ END DEBUG ############*/
test_input[33288:33295] = '{32'hc29de789, 32'h42a01c01, 32'h421ef8cd, 32'hc1e2a707, 32'hc11930bf, 32'hc2914dea, 32'hc1e4f7f3, 32'hc0c7f303};
test_label[4161] = '{32'hc0c7f303};
test_output[4161] = '{32'h42ac9b31};
/*############ DEBUG ############
test_input[33288:33295] = '{-78.952218329, 80.0546925131, 39.7429695246, -28.3315563035, -9.5744009439, -72.6521785082, -28.6210682887, -6.2484147464};
test_label[4161] = '{-6.2484147464};
test_output[4161] = '{86.3031072595};
############ END DEBUG ############*/
test_input[33296:33303] = '{32'h4254f34f, 32'h403aad68, 32'hc27fcf71, 32'hc29983a9, 32'hc086c994, 32'h42c142cc, 32'hc20504a5, 32'h41c2975f};
test_label[4162] = '{32'h41c2975f};
test_output[4162] = '{32'h42909cf4};
/*############ DEBUG ############
test_input[33296:33303] = '{53.2376061678, 2.91683387724, -63.9525796192, -76.7571481845, -4.21210663809, 96.6304639808, -33.2545374759, 24.323912385};
test_label[4162] = '{24.323912385};
test_output[4162] = '{72.3065515958};
############ END DEBUG ############*/
test_input[33304:33311] = '{32'hc2424c3f, 32'hc1e32e79, 32'hc227de9a, 32'hc11d0bc1, 32'hc26ecc85, 32'hc0e10cf4, 32'hc1c25641, 32'h411459b0};
test_label[4163] = '{32'hc0e10cf4};
test_output[4163] = '{32'h41827015};
/*############ DEBUG ############
test_input[33304:33311] = '{-48.5744593889, -28.3976923698, -41.9673830677, -9.81536944412, -59.6997265728, -7.03283111618, -24.292117089, 9.2718965981};
test_label[4163] = '{-7.03283111618};
test_output[4163] = '{16.3047278024};
############ END DEBUG ############*/
test_input[33312:33319] = '{32'hc126fb0c, 32'hc24e0507, 32'hc2a5c509, 32'hc124b8d1, 32'h429108e2, 32'hc20cbfa6, 32'h413f5007, 32'hc284d982};
test_label[4164] = '{32'hc20cbfa6};
test_output[4164] = '{32'h42d768b5};
/*############ DEBUG ############
test_input[33312:33319] = '{-10.436290722, -51.5049095061, -82.8848336374, -10.2951211215, 72.5173486347, -35.1871575179, 11.9570378223, -66.424820137};
test_label[4164] = '{-35.1871575179};
test_output[4164] = '{107.704506153};
############ END DEBUG ############*/
test_input[33320:33327] = '{32'h428aa6b0, 32'hc259062d, 32'h415b1484, 32'hc2a1e4ee, 32'hc2ad08d1, 32'hc19be4ff, 32'h4213e149, 32'hc21d6fa2};
test_label[4165] = '{32'h428aa6b0};
test_output[4165] = '{32'h281e0000};
/*############ DEBUG ############
test_input[33320:33327] = '{69.3255639675, -54.2560318941, 13.6925086048, -80.9471320746, -86.5172219507, -19.4868150734, 36.9700060967, -39.3590156957};
test_label[4165] = '{69.3255639675};
test_output[4165] = '{8.77076189454e-15};
############ END DEBUG ############*/
test_input[33328:33335] = '{32'hc187f8ea, 32'h420d5ee2, 32'hc2a7b3f2, 32'h4197b621, 32'hc20f669b, 32'h4274ff51, 32'h42896e95, 32'hc2aaeea5};
test_label[4166] = '{32'hc2aaeea5};
test_output[4166] = '{32'h431a2ec3};
/*############ DEBUG ############
test_input[33328:33335] = '{-16.9965394768, 35.3426604571, -83.8514531713, 18.9639302137, -35.8501998497, 61.2493312163, 68.7159799636, -85.4661041691};
test_label[4166] = '{-85.4661041691};
test_output[4166] = '{154.182655811};
############ END DEBUG ############*/
test_input[33336:33343] = '{32'h42c6b43a, 32'h423150f7, 32'hc2a2d686, 32'hc28ea482, 32'h426575ac, 32'h41ab1a65, 32'hc1412df1, 32'h41c82512};
test_label[4167] = '{32'h41ab1a65};
test_output[4167] = '{32'h429beda0};
/*############ DEBUG ############
test_input[33336:33343] = '{99.3520014312, 44.32906709, -81.4189886735, -71.3213025882, 57.3649143083, 21.3878886414, -12.0737163013, 25.0181002518};
test_label[4167] = '{21.3878886414};
test_output[4167] = '{77.9641127898};
############ END DEBUG ############*/
test_input[33344:33351] = '{32'h422ffd68, 32'h428161d6, 32'hc2bcc7cc, 32'hc2b0de41, 32'h4221fda9, 32'hc1a51aeb, 32'hc2107875, 32'hc2241f09};
test_label[4168] = '{32'h4221fda9};
test_output[4168] = '{32'h41c18c04};
/*############ DEBUG ############
test_input[33344:33351] = '{43.9974676502, 64.6910833262, -94.390226479, -88.4340924124, 40.4977161004, -20.6381427794, -36.1176351677, -41.0303066913};
test_label[4168] = '{40.4977161004};
test_output[4168] = '{24.1933672269};
############ END DEBUG ############*/
test_input[33352:33359] = '{32'h41f7993e, 32'h42b4ea7e, 32'h4255f612, 32'h4298a9b1, 32'hc2b6bfe4, 32'h4213a15d, 32'h42c5d86f, 32'hc2c62b7e};
test_label[4169] = '{32'h41f7993e};
test_output[4169] = '{32'h4287f23b};
/*############ DEBUG ############
test_input[33352:33359] = '{30.9498260856, 90.4579914351, 53.4903021119, 76.3314287692, -91.3747897376, 36.9075814601, 98.9227248907, -99.0849422176};
test_label[4169] = '{30.9498260856};
test_output[4169] = '{67.9731095552};
############ END DEBUG ############*/
test_input[33360:33367] = '{32'h42bf7f4c, 32'hc20aade9, 32'h42591174, 32'hc2880216, 32'h4218c8ef, 32'hc2585650, 32'hc1dcbcf4, 32'hc28325ae};
test_label[4170] = '{32'h4218c8ef};
test_output[4170] = '{32'h426635a9};
/*############ DEBUG ############
test_input[33360:33367] = '{95.7486289869, -34.6698345162, 54.2670458081, -68.004073204, 38.1962245845, -54.0842906371, -27.592261466, -65.5735954042};
test_label[4170] = '{38.1962245845};
test_output[4170] = '{57.5524044025};
############ END DEBUG ############*/
test_input[33368:33375] = '{32'hc1a850fb, 32'h41aa51c2, 32'hc1f789eb, 32'h426c3014, 32'h41a286ec, 32'h40d46390, 32'h4286ea29, 32'hc205d060};
test_label[4171] = '{32'h40d46390};
test_output[4171] = '{32'h4273481b};
/*############ DEBUG ############
test_input[33368:33375] = '{-21.0395407388, 21.2899201211, -30.942342128, 59.0469496275, 20.315880157, 6.63715370912, 67.4573466485, -33.4534929082};
test_label[4171] = '{6.63715370912};
test_output[4171] = '{60.8204154561};
############ END DEBUG ############*/
test_input[33376:33383] = '{32'hc139a874, 32'hc28e51ac, 32'hc25cb5c7, 32'hc2be8fd8, 32'h4298ee77, 32'hc261fd74, 32'hc1a578ea, 32'h41d074dd};
test_label[4172] = '{32'h4298ee77};
test_output[4172] = '{32'h80000000};
/*############ DEBUG ############
test_input[33376:33383] = '{-11.6036265659, -71.1595160126, -55.1775180066, -95.2809413082, 76.4657481933, -56.4975112103, -20.6840392744, 26.0570629279};
test_label[4172] = '{76.4657481933};
test_output[4172] = '{-0.0};
############ END DEBUG ############*/
test_input[33384:33391] = '{32'hc083cadb, 32'h42108b64, 32'hc29ec619, 32'h423ed5b5, 32'h42abf410, 32'hc259dc6f, 32'h4109eb49, 32'h4299067a};
test_label[4173] = '{32'hc083cadb};
test_output[4173] = '{32'h42b430c8};
/*############ DEBUG ############
test_input[33384:33391] = '{-4.11851263674, 36.136124082, -79.3869097613, 47.7086966065, 85.9766862737, -54.4652684825, 8.61994238437, 76.512651651};
test_label[4173] = '{-4.11851263674};
test_output[4173] = '{90.0952765003};
############ END DEBUG ############*/
test_input[33392:33399] = '{32'h41f4925e, 32'h41cfaf9d, 32'h42187e5c, 32'hc292e7eb, 32'hc293e764, 32'h4214812e, 32'h40e6cd4c, 32'hc2966156};
test_label[4174] = '{32'h42187e5c};
test_output[4174] = '{32'h3ea0f7d6};
/*############ DEBUG ############
test_input[33392:33399] = '{30.5714679481, 25.9607493164, 38.1233972802, -73.4529628097, -73.9519324223, 37.1261527682, 7.21256066307, -75.1901116461};
test_label[4174] = '{38.1233972802};
test_output[4174] = '{0.314390830119};
############ END DEBUG ############*/
test_input[33400:33407] = '{32'h429fc47e, 32'h428e9a47, 32'hc25e5bf7, 32'h424c44dd, 32'hc25ec733, 32'h40df293b, 32'h429b69ff, 32'h42a5b811};
test_label[4175] = '{32'h424c44dd};
test_output[4175] = '{32'h41fec7b0};
/*############ DEBUG ############
test_input[33400:33407] = '{79.8837734973, 71.3013222453, -55.5898109598, 51.067250175, -55.6945314859, 6.97378310973, 77.7070230911, 82.8595033149};
test_label[4175] = '{51.067250175};
test_output[4175] = '{31.8475031453};
############ END DEBUG ############*/
test_input[33408:33415] = '{32'hc2b53e5f, 32'h42bbc8e4, 32'h4283b161, 32'h42b53925, 32'hc254a91a, 32'h4289795b, 32'h4269c2f6, 32'hc28bbfdd};
test_label[4176] = '{32'h4289795b};
test_output[4176] = '{32'h41c989b8};
/*############ DEBUG ############
test_input[33408:33415] = '{-90.6218223409, 93.8923610763, 65.8464421858, 90.6116083231, -53.1651382341, 68.7370252128, 58.4403901551, -69.8747339849};
test_label[4176] = '{68.7370252128};
test_output[4176] = '{25.1922461623};
############ END DEBUG ############*/
test_input[33416:33423] = '{32'hc27b0df0, 32'h42bfa452, 32'hc2c16043, 32'hc203f02e, 32'h415c4dad, 32'hc2a03c94, 32'h41e0c209, 32'hc2490b4c};
test_label[4177] = '{32'hc2c16043};
test_output[4177] = '{32'h4340824b};
/*############ DEBUG ############
test_input[33416:33423] = '{-62.7636101, 95.820941545, -96.6880124872, -32.9845492334, 13.7689634145, -80.1183196845, 28.0947438387, -50.2610333501};
test_label[4177] = '{-96.6880124872};
test_output[4177] = '{192.508954032};
############ END DEBUG ############*/
test_input[33424:33431] = '{32'hc24ec3ae, 32'hc20dd8ae, 32'hc23a9469, 32'h419eadba, 32'h42389e23, 32'hc2c56aef, 32'h4198ccf3, 32'h4289e771};
test_label[4178] = '{32'hc24ec3ae};
test_output[4178] = '{32'h42f14948};
/*############ DEBUG ############
test_input[33424:33431] = '{-51.6910919051, -35.4616025151, -46.6449303556, 19.8348274853, 46.1544308226, -98.7088564499, 19.1000729089, 68.9520371575};
test_label[4178] = '{-51.6910919051};
test_output[4178] = '{120.643129063};
############ END DEBUG ############*/
test_input[33432:33439] = '{32'hc27943db, 32'hc22c76ed, 32'h429d61d7, 32'hc0a78dae, 32'hc2b2291f, 32'hc1bbc6b3, 32'hc2b31092, 32'hc2b99e96};
test_label[4179] = '{32'hc22c76ed};
test_output[4179] = '{32'h42f39d4e};
/*############ DEBUG ############
test_input[33432:33439] = '{-62.3162638988, -43.1161400568, 78.691094217, -5.23604498494, -89.080312241, -23.4720206719, -89.5323620646, -92.8097344373};
test_label[4179] = '{-43.1161400568};
test_output[4179] = '{121.807234274};
############ END DEBUG ############*/
test_input[33440:33447] = '{32'h429e7b78, 32'h42c0a448, 32'hc2a1889b, 32'h4274ecb1, 32'h4221a601, 32'hc2a07a0d, 32'hc20f37af, 32'hc29ae8b8};
test_label[4180] = '{32'h4274ecb1};
test_output[4180] = '{32'h420c5be0};
/*############ DEBUG ############
test_input[33440:33447] = '{79.2411512115, 96.3208653435, -80.7668079272, 61.2311438551, 40.4121145846, -80.2383828889, -35.8043798981, -77.454528198};
test_label[4180] = '{61.2311438551};
test_output[4180] = '{35.0897215266};
############ END DEBUG ############*/
test_input[33448:33455] = '{32'h400da771, 32'h42854928, 32'hc29af689, 32'h41b111f1, 32'hc2457c93, 32'hc21bfc00, 32'hc1e6207d, 32'h4247744f};
test_label[4181] = '{32'hc21bfc00};
test_output[4181] = '{32'h42d34728};
/*############ DEBUG ############
test_input[33448:33455] = '{2.21334489811, 66.6428845094, -77.4815167205, 22.1337606561, -49.3716552713, -38.9960948572, -28.7658639386, 49.8635844327};
test_label[4181] = '{-38.9960948572};
test_output[4181] = '{105.638979418};
############ END DEBUG ############*/
test_input[33456:33463] = '{32'hc2c48caf, 32'h42580186, 32'h42024cae, 32'hc2522cbb, 32'h42a0a4fa, 32'h42b90187, 32'h420fa43d, 32'hc267f249};
test_label[4182] = '{32'hc2c48caf};
test_output[4182] = '{32'h433ec71c};
/*############ DEBUG ############
test_input[33456:33463] = '{-98.2747755386, 54.0014892524, 32.5748816063, -52.5436823552, 80.3222227904, 92.5029847035, 35.9103907359, -57.9866084282};
test_label[4182] = '{-98.2747755386};
test_output[4182] = '{190.77776537};
############ END DEBUG ############*/
test_input[33464:33471] = '{32'hc2c3d225, 32'h428168d7, 32'hc1816b2e, 32'hc28785c7, 32'h4138a884, 32'h4288b63c, 32'h42479517, 32'hc2136168};
test_label[4183] = '{32'h428168d7};
test_output[4183] = '{32'h406b5094};
/*############ DEBUG ############
test_input[33464:33471] = '{-97.9104365443, 64.7047637327, -16.1773334298, -67.7612829028, 11.5411413027, 68.3559271233, 49.8955952504, -36.845123719};
test_label[4183] = '{64.7047637327};
test_output[4183] = '{3.6767930451};
############ END DEBUG ############*/
test_input[33472:33479] = '{32'hc29feb78, 32'hc21ad04a, 32'hc2b59697, 32'hc2a6e86e, 32'h421e7570, 32'hc21a6765, 32'hc2503609, 32'hc213fd8e};
test_label[4184] = '{32'h421e7570};
test_output[4184] = '{32'h80000000};
/*############ DEBUG ############
test_input[33472:33479] = '{-79.9598997839, -38.7034079841, -90.794121696, -83.4539632982, 39.6146856783, -38.6009699871, -52.0527673975, -36.9976117402};
test_label[4184] = '{39.6146856783};
test_output[4184] = '{-0.0};
############ END DEBUG ############*/
test_input[33480:33487] = '{32'h41c5fa9c, 32'h42298c5b, 32'h4192b383, 32'h42024dc5, 32'hc29a8f0d, 32'hc278dd31, 32'h4138483b, 32'hc2c72d68};
test_label[4185] = '{32'hc2c72d68};
test_output[4185] = '{32'h430df9ce};
/*############ DEBUG ############
test_input[33480:33487] = '{24.7473669297, 42.3870665678, 18.337652906, 32.5759474839, -77.2793990892, -62.216005538, 11.5176342565, -99.5886814466};
test_label[4185] = '{-99.5886814466};
test_output[4185] = '{141.975802873};
############ END DEBUG ############*/
test_input[33488:33495] = '{32'hc040b48a, 32'hc2be1602, 32'h42c3049a, 32'h42bc0fc6, 32'hc2bff20f, 32'h41ec17e0, 32'h426ae485, 32'hc283335a};
test_label[4186] = '{32'hc2be1602};
test_output[4186] = '{32'h43409516};
/*############ DEBUG ############
test_input[33488:33495] = '{-3.01101914958, -95.0429856492, 97.5089907989, 94.0308038208, -95.9727734662, 29.5116576718, 58.7231649369, -65.6002933955};
test_label[4186] = '{-95.0429856492};
test_output[4186] = '{192.58237307};
############ END DEBUG ############*/
test_input[33496:33503] = '{32'hc226a195, 32'h41ab11ae, 32'hc2864142, 32'h42b28221, 32'h42c644ea, 32'hc2bc6e62, 32'h41cdd0c7, 32'h41bd8b2a};
test_label[4187] = '{32'hc2864142};
test_output[4187] = '{32'h43264319};
/*############ DEBUG ############
test_input[33496:33503] = '{-41.6577946654, 21.3836320854, -67.1274549441, 89.2541615369, 99.1345967035, -94.2155877266, 25.7269415338, 23.6929520028};
test_label[4187] = '{-67.1274549441};
test_output[4187] = '{166.262102812};
############ END DEBUG ############*/
test_input[33504:33511] = '{32'hc2857be7, 32'hc2c7f39c, 32'hc25843f8, 32'h417460bf, 32'hc24194aa, 32'hc177173a, 32'h42633228, 32'hc1e38bd0};
test_label[4188] = '{32'hc2c7f39c};
test_output[4188] = '{32'h431cc658};
/*############ DEBUG ############
test_input[33504:33511] = '{-66.7419960749, -99.9757982096, -54.0663761835, 15.2736195735, -48.3951802479, -15.4431705686, 56.798979497, -28.4432670043};
test_label[4188] = '{-99.9757982096};
test_output[4188] = '{156.774777707};
############ END DEBUG ############*/
test_input[33512:33519] = '{32'hc18b4265, 32'h425a38a1, 32'h42b9fd6d, 32'hc1d8c529, 32'hc2b7d737, 32'h42b6581e, 32'hc155134a, 32'hc2844d03};
test_label[4189] = '{32'hc1d8c529};
test_output[4189] = '{32'h42f07b65};
/*############ DEBUG ############
test_input[33512:33519] = '{-17.4074200119, 54.5553004231, 92.9949730493, -27.0962692974, -91.9203384784, 91.1721024193, -13.3172088881, -66.1504151351};
test_label[4189] = '{-27.0962692974};
test_output[4189] = '{120.241007397};
############ END DEBUG ############*/
test_input[33520:33527] = '{32'hc09dc884, 32'h421e5b30, 32'hc2949869, 32'h425e19bd, 32'h41618316, 32'h4230e78c, 32'h4279f4cf, 32'h4211cb3c};
test_label[4190] = '{32'h41618316};
test_output[4190] = '{32'h42419502};
/*############ DEBUG ############
test_input[33520:33527] = '{-4.93072701259, 39.5890518951, -74.297674684, 55.5251352787, 14.0945032818, 44.2261214693, 62.4890725677, 36.4484708576};
test_label[4190] = '{14.0945032818};
test_output[4190] = '{48.3955142181};
############ END DEBUG ############*/
test_input[33528:33535] = '{32'h425b838c, 32'hc25c0255, 32'hc2b2b8b2, 32'hc29f7a8d, 32'hc20dd93d, 32'h4051ce5f, 32'h424fc5c1, 32'hc117500a};
test_label[4191] = '{32'hc20dd93d};
test_output[4191] = '{32'h42b4c8e4};
/*############ DEBUG ############
test_input[33528:33535] = '{54.8784654509, -55.0022766768, -89.3607307931, -79.7393537885, -35.4621471259, 3.27822080174, 51.9431185869, -9.45704049107};
test_label[4191] = '{-35.4621471259};
test_output[4191] = '{90.3923624456};
############ END DEBUG ############*/
test_input[33536:33543] = '{32'h42a465af, 32'h40bc47d7, 32'h4120305b, 32'h41431603, 32'hc2ad3738, 32'h42b2a254, 32'hc281abfc, 32'hc2160d5c};
test_label[4192] = '{32'hc2160d5c};
test_output[4192] = '{32'h42fda96c};
/*############ DEBUG ############
test_input[33536:33543] = '{82.1986018237, 5.88376968412, 10.0118054512, 12.192873745, -86.6078483462, 89.3170483345, -64.8359062562, -37.5130458344};
test_label[4192] = '{-37.5130458344};
test_output[4192] = '{126.830903865};
############ END DEBUG ############*/
test_input[33544:33551] = '{32'hc2409186, 32'h42c1009d, 32'h42152542, 32'hc292bbc5, 32'hc2c013b4, 32'hc2ac6e1b, 32'hc2955061, 32'hc2c4b8e4};
test_label[4193] = '{32'hc2c4b8e4};
test_output[4193] = '{32'h4342dcc0};
/*############ DEBUG ############
test_input[33544:33551] = '{-48.142112356, 96.5011983427, 37.2863827327, -73.3667370492, -96.0384810907, -86.215047625, -74.6569862378, -98.3611134982};
test_label[4193] = '{-98.3611134982};
test_output[4193] = '{194.862311841};
############ END DEBUG ############*/
test_input[33552:33559] = '{32'h42ab099d, 32'h41b31ff2, 32'hc046d1b1, 32'hc1f28399, 32'hc1552e9e, 32'hc27f4c7f, 32'hc1b6aef1, 32'hc2491f92};
test_label[4194] = '{32'hc2491f92};
test_output[4194] = '{32'h4307ccb3};
/*############ DEBUG ############
test_input[33552:33559] = '{85.5187725787, 22.3905974987, -3.1065485438, -30.3142558648, -13.3238815111, -63.8247014457, -22.8354215356, -50.2808310279};
test_label[4194] = '{-50.2808310279};
test_output[4194] = '{135.799603607};
############ END DEBUG ############*/
test_input[33560:33567] = '{32'h40d1be36, 32'hc29870ea, 32'h4244fdfb, 32'hc29f44d6, 32'hc28f884d, 32'hc29b6e23, 32'h3f6bcf60, 32'h428218cc};
test_label[4195] = '{32'hc29b6e23};
test_output[4195] = '{32'h430ec377};
/*############ DEBUG ############
test_input[33560:33567] = '{6.55446891818, -76.2205316439, 49.2480295844, -79.6344465141, -71.7662092197, -77.7151099521, 0.921133019114, 65.0484313351};
test_label[4195] = '{-77.7151099521};
test_output[4195] = '{142.763541425};
############ END DEBUG ############*/
test_input[33568:33575] = '{32'h42700d37, 32'h42adab39, 32'hc0b12585, 32'hc1185cbb, 32'hc2bf62e5, 32'h422ec72b, 32'hc1b8831b, 32'hc20e71fa};
test_label[4196] = '{32'hc0b12585};
test_output[4196] = '{32'h42b8bd92};
/*############ DEBUG ############
test_input[33568:33575] = '{60.0129066206, 86.8344205421, -5.53583022175, -9.52263968972, -95.6931537255, 43.6944995058, -23.0640159617, -35.6113045053};
test_label[4196] = '{-5.53583022175};
test_output[4196] = '{92.3702507639};
############ END DEBUG ############*/
test_input[33576:33583] = '{32'h42af19ab, 32'h415056f9, 32'hc2be528f, 32'hc264b5ed, 32'hc290ac10, 32'h425dc891, 32'h4254a0bf, 32'h42a84ad3};
test_label[4197] = '{32'h425dc891};
test_output[4197] = '{32'h42008c40};
/*############ DEBUG ############
test_input[33576:33583] = '{87.5501289516, 13.0212334428, -95.1612469119, -57.1776615572, -72.336059973, 55.4458652525, 53.1569797139, 84.1461397689};
test_label[4197] = '{55.4458652525};
test_output[4197] = '{32.1369635854};
############ END DEBUG ############*/
test_input[33584:33591] = '{32'h422e2fb9, 32'hc2a68c33, 32'h429249b6, 32'hc260df07, 32'hc2a6a942, 32'hc23fd2fc, 32'hc1005c3f, 32'hc2c6bfb3};
test_label[4198] = '{32'h422e2fb9};
test_output[4198] = '{32'h41ecc766};
/*############ DEBUG ############
test_input[33584:33591] = '{43.5466023667, -83.2738266087, 73.1439657542, -56.2177995459, -83.3305782039, -47.9560410967, -8.02252137309, -99.3744118896};
test_label[4198] = '{43.5466023667};
test_output[4198] = '{29.5973633875};
############ END DEBUG ############*/
test_input[33592:33599] = '{32'h3f7cbe62, 32'h429eee63, 32'hc208a1dd, 32'hc2be93ac, 32'hc1664bad, 32'h40d32b35, 32'h42c445af, 32'hc2c02bc4};
test_label[4199] = '{32'hc2be93ac};
test_output[4199] = '{32'h43416cae};
/*############ DEBUG ############
test_input[33592:33599] = '{0.987280023289, 79.4656013018, -34.1580705693, -95.2884248034, -14.3934752124, 6.59902446532, 98.1361032983, -96.0854828271};
test_label[4199] = '{-95.2884248034};
test_output[4199] = '{193.424528109};
############ END DEBUG ############*/
test_input[33600:33607] = '{32'hc2873b92, 32'hc1b7663c, 32'hc248b08f, 32'h42c0fe30, 32'hc2b71bfb, 32'h426d4455, 32'hc290dd24, 32'hc29c4a7a};
test_label[4200] = '{32'hc1b7663c};
test_output[4200] = '{32'h42eed7bf};
/*############ DEBUG ############
test_input[33600:33607] = '{-67.6163466734, -22.9249185598, -50.1724198424, 96.4964585858, -91.5546528778, 59.3167303565, -72.4319144792, -78.1454582315};
test_label[4200] = '{-22.9249185598};
test_output[4200] = '{119.421377146};
############ END DEBUG ############*/
test_input[33608:33615] = '{32'hc213a3ca, 32'hc2386b67, 32'h42c10105, 32'h420b3eb3, 32'hc21adb34, 32'h424e5a9f, 32'h428ffcf7, 32'hc1a2dce2};
test_label[4201] = '{32'h424e5a9f};
test_output[4201] = '{32'h4233a76c};
/*############ DEBUG ############
test_input[33608:33615] = '{-36.9099508901, -46.1048860057, 96.5019939593, 34.8112279863, -38.7140640408, 51.5884965756, 71.9940703712, -20.3578524782};
test_label[4201] = '{51.5884965756};
test_output[4201] = '{44.9134973838};
############ END DEBUG ############*/
test_input[33616:33623] = '{32'h4221d638, 32'h41bdd4de, 32'h4230a259, 32'hc27f60a8, 32'h4180fe79, 32'h41b104c7, 32'hc291233e, 32'hc28a1c95};
test_label[4202] = '{32'hc28a1c95};
test_output[4202] = '{32'h42e27a44};
/*############ DEBUG ############
test_input[33616:33623] = '{40.4591984718, 23.7289395454, 44.1585426961, -63.8443925807, 16.124254947, 22.1273332658, -72.5688351902, -69.0558223839};
test_label[4202] = '{-69.0558223839};
test_output[4202] = '{113.238803754};
############ END DEBUG ############*/
test_input[33624:33631] = '{32'h42919dd5, 32'h412c280a, 32'hc2a7938f, 32'hc1e1e9e6, 32'h409c0cae, 32'h42876bad, 32'hc2823b7a, 32'h42b2150c};
test_label[4203] = '{32'h42919dd5};
test_output[4203] = '{32'h4181dcdb};
/*############ DEBUG ############
test_input[33624:33631] = '{72.8082688985, 10.7597749633, -83.7882026118, -28.2392080637, 4.87654777085, 67.7103008536, -65.1161657049, 89.0411081084};
test_label[4203] = '{72.8082688985};
test_output[4203] = '{16.2328392995};
############ END DEBUG ############*/
test_input[33632:33639] = '{32'hc2ab86c6, 32'h41e57b8c, 32'h417673bd, 32'hc1e38f0d, 32'h42b63d4a, 32'hc1299b55, 32'h41718f4a, 32'h4252b5e8};
test_label[4204] = '{32'h417673bd};
test_output[4204] = '{32'h42976ed2};
/*############ DEBUG ############
test_input[33632:33639] = '{-85.7632290625, 28.6853264617, 15.4032567204, -28.444849456, 91.1197053829, -10.6004229657, 15.0974823922, 52.6776416017};
test_label[4204] = '{15.4032567204};
test_output[4204] = '{75.7164486625};
############ END DEBUG ############*/
test_input[33640:33647] = '{32'hc190a640, 32'hc2a9f83d, 32'hc1db3198, 32'hc1aaed58, 32'h4281b0fd, 32'h42afee83, 32'h423b9e36, 32'hc2368b5d};
test_label[4205] = '{32'hc190a640};
test_output[4205] = '{32'h42d41813};
/*############ DEBUG ############
test_input[33640:33647] = '{-18.0811769927, -84.9848436111, -27.399215066, -21.3658900381, 64.8456835959, 87.9658412002, 46.9045041651, -45.6360954593};
test_label[4205] = '{-18.0811769927};
test_output[4205] = '{106.047018193};
############ END DEBUG ############*/
test_input[33648:33655] = '{32'h420b63d8, 32'hc27225d6, 32'hc1e7fd0e, 32'hc184230b, 32'hc26870f8, 32'hc2146c70, 32'h42343bbd, 32'h42ae2114};
test_label[4206] = '{32'hc184230b};
test_output[4206] = '{32'h42cf29d7};
/*############ DEBUG ############
test_input[33648:33655] = '{34.8475042389, -60.5369505139, -28.9985618238, -16.5171107565, -58.1103224419, -37.1058974256, 45.0583376738, 87.0646059281};
test_label[4206] = '{-16.5171107565};
test_output[4206] = '{103.581716685};
############ END DEBUG ############*/
test_input[33656:33663] = '{32'hc22ca4ee, 32'hc29805a6, 32'hc18474f6, 32'h4229abd7, 32'h424f40e8, 32'h4240cb12, 32'hc2283caa, 32'hc2c72a7c};
test_label[4207] = '{32'h4229abd7};
test_output[4207] = '{32'h4116c164};
/*############ DEBUG ############
test_input[33656:33663] = '{-43.1610640153, -76.0110295831, -16.5571094665, 42.4178119357, 51.8133861902, 48.1983099621, -42.0592407102, -99.5829754627};
test_label[4207] = '{42.4178119357};
test_output[4207] = '{9.4222142034};
############ END DEBUG ############*/
test_input[33664:33671] = '{32'h42361983, 32'hc1b8249d, 32'hc14f1b63, 32'hc29f128f, 32'hc109bf3c, 32'h42bb228f, 32'hc2052a97, 32'h423595c7};
test_label[4208] = '{32'hc29f128f};
test_output[4208] = '{32'h432d1a8f};
/*############ DEBUG ############
test_input[33664:33671] = '{45.5249123544, -23.0178780099, -12.9441859244, -79.5362465749, -8.60918851841, 93.5674959357, -33.2915925108, 45.3962675082};
test_label[4208] = '{-79.5362465749};
test_output[4208] = '{173.103742511};
############ END DEBUG ############*/
test_input[33672:33679] = '{32'h42427c03, 32'h42a8fab3, 32'hc24e1c06, 32'h41bbfcc6, 32'hc2a92a33, 32'hc2391b23, 32'hc29549cb, 32'hc28945ec};
test_label[4209] = '{32'hc2a92a33};
test_output[4209] = '{32'h43291273};
/*############ DEBUG ############
test_input[33672:33679] = '{48.621103898, 84.4896497392, -51.5273668453, 23.4984242441, -84.5824227944, -46.2765019935, -74.6441247724, -68.6365684557};
test_label[4209] = '{-84.5824227944};
test_output[4209] = '{169.072072534};
############ END DEBUG ############*/
test_input[33680:33687] = '{32'h42565fbb, 32'h41bce9ac, 32'h41abda6b, 32'hc2c078e9, 32'h40d20a8b, 32'hc067fcd3, 32'hc24d02a1, 32'h42add197};
test_label[4210] = '{32'h41bce9ac};
test_output[4210] = '{32'h427d2e58};
/*############ DEBUG ############
test_input[33680:33687] = '{53.5934853193, 23.6140976567, 21.4816502536, -96.2361559935, 6.56378712721, -3.62480615105, -51.2525658546, 86.9093560043};
test_label[4210] = '{23.6140976567};
test_output[4210] = '{63.2952583476};
############ END DEBUG ############*/
test_input[33688:33695] = '{32'h4254f53b, 32'h42a196cd, 32'h41faa1c1, 32'h42456162, 32'h42244f63, 32'h429fd0be, 32'hc0c00e38, 32'h41413ce4};
test_label[4211] = '{32'h4254f53b};
test_output[4211] = '{32'h41df3341};
/*############ DEBUG ############
test_input[33688:33695] = '{53.2394835071, 80.7945298905, 31.3289822495, 49.3451022919, 41.0775263028, 79.9077027983, -6.00173582369, 12.0773659326};
test_label[4211] = '{53.2394835071};
test_output[4211] = '{27.9000257564};
############ END DEBUG ############*/
test_input[33696:33703] = '{32'h42214065, 32'hc20b986e, 32'hc18d03d2, 32'hc2c7c5b6, 32'h413e0713, 32'h425fbd2c, 32'h40a1663d, 32'hc20592fc};
test_label[4212] = '{32'h413e0713};
test_output[4212] = '{32'h42303b68};
/*############ DEBUG ############
test_input[33696:33703] = '{40.3128870117, -34.8988573582, -17.6268663272, -99.8861526031, 11.8767275709, 55.9347395848, 5.04373038812, -33.3935389538};
test_label[4212] = '{11.8767275709};
test_output[4212] = '{44.0580121781};
############ END DEBUG ############*/
test_input[33704:33711] = '{32'hc2b6c1f2, 32'hbfaf7485, 32'h4143b75e, 32'h42842dd3, 32'h428344d5, 32'h4242ec52, 32'hc23a776b, 32'h42b3c6dd};
test_label[4213] = '{32'h4242ec52};
test_output[4213] = '{32'h4224a168};
/*############ DEBUG ############
test_input[33704:33711] = '{-91.3787968262, -1.37074340195, 12.2322669874, 66.0895025426, 65.6344378548, 48.7307825115, -46.6166193574, 89.8884054598};
test_label[4213] = '{48.7307825115};
test_output[4213] = '{41.1576229484};
############ END DEBUG ############*/
test_input[33712:33719] = '{32'hc293562f, 32'hc171483d, 32'hc2b53f44, 32'h42c5ffc8, 32'h428ed3ca, 32'hc23ededc, 32'hc28490bd, 32'hc2a41f89};
test_label[4214] = '{32'hc171483d};
test_output[4214] = '{32'h42e428cf};
/*############ DEBUG ############
test_input[33712:33719] = '{-73.6683268318, -15.0801361149, -90.623566783, 98.9995708154, 71.4136535392, -47.7176361408, -66.2826927263, -82.0615910984};
test_label[4214] = '{-15.0801361149};
test_output[4214] = '{114.07970693};
############ END DEBUG ############*/
test_input[33720:33727] = '{32'h42be8199, 32'h42a1c9fa, 32'h429a9322, 32'h420d9316, 32'h41b00473, 32'h4252924e, 32'hc2ad7204, 32'hc28b3420};
test_label[4215] = '{32'h420d9316};
test_output[4215] = '{32'h426f701d};
/*############ DEBUG ############
test_input[33720:33727] = '{95.2531214708, 80.8944839806, 77.2873668826, 35.3936371398, 22.002172307, 52.6428756633, -86.7226901186, -69.6018077299};
test_label[4215] = '{35.3936371398};
test_output[4215] = '{59.8594849276};
############ END DEBUG ############*/
test_input[33728:33735] = '{32'h41cc04e7, 32'h41f63c5e, 32'h421d40ce, 32'h40aff599, 32'hc1d15098, 32'h42b76987, 32'hc2ae6f81, 32'hc22687b9};
test_label[4216] = '{32'h41f63c5e};
test_output[4216] = '{32'h4273b4df};
/*############ DEBUG ############
test_input[33728:33735] = '{25.5023940669, 30.7794762716, 39.3132846679, 5.49872994872, -26.164353106, 91.7061078538, -87.2177781698, -41.632540232};
test_label[4216] = '{30.7794762716};
test_output[4216] = '{60.9266315822};
############ END DEBUG ############*/
test_input[33736:33743] = '{32'hc2a20426, 32'hc20b8acb, 32'h42bbb179, 32'hc2648758, 32'hc2541179, 32'h4205e031, 32'h4281cf67, 32'h41f59602};
test_label[4217] = '{32'h4281cf67};
test_output[4217] = '{32'h41e78846};
/*############ DEBUG ############
test_input[33736:33743] = '{-81.0081037703, -34.8855396538, 93.8466252906, -57.1321703949, -53.0170638734, 33.4689387792, 64.90508466, 30.6982466296};
test_label[4217] = '{64.90508466};
test_output[4217] = '{28.9415406305};
############ END DEBUG ############*/
test_input[33744:33751] = '{32'hc231c5c9, 32'hc2146775, 32'hc189af1f, 32'h42a640e9, 32'hc18766dd, 32'hc2121857, 32'hc26b13fb, 32'hc2ab796f};
test_label[4218] = '{32'hc2ab796f};
test_output[4218] = '{32'h4328dd2c};
/*############ DEBUG ############
test_input[33744:33751] = '{-44.4431494919, -37.1010326112, -17.2105086981, 83.1267754275, -16.9252252842, -36.5237691114, -58.7695140683, -85.737173092};
test_label[4218] = '{-85.737173092};
test_output[4218] = '{168.863948519};
############ END DEBUG ############*/
test_input[33752:33759] = '{32'h42059a7e, 32'hc28e09bc, 32'h4287a3ff, 32'hc130efa0, 32'h41f6b8d3, 32'hc22e2061, 32'hc2471225, 32'hc2b03b51};
test_label[4219] = '{32'hc2b03b51};
test_output[4219] = '{32'h431befa8};
/*############ DEBUG ############
test_input[33752:33759] = '{33.4008704628, -71.0190103584, 67.8203077998, -11.0585024147, 30.8402458361, -43.5316195788, -49.7677187951, -88.1158551147};
test_label[4219] = '{-88.1158551147};
test_output[4219] = '{155.936162914};
############ END DEBUG ############*/
test_input[33760:33767] = '{32'h429a0e77, 32'hc2aa6dd5, 32'hc2306250, 32'h4296d14d, 32'hbf8633de, 32'hc19b89f8, 32'h3f91539f, 32'h414dae43};
test_label[4220] = '{32'hc19b89f8};
test_output[4220] = '{32'h42c14d74};
/*############ DEBUG ############
test_input[33760:33767] = '{77.0282515077, -85.2145149008, -44.096008139, 75.4087897663, -1.0484578412, -19.4423682196, 1.1353644488, 12.855044055};
test_label[4220] = '{-19.4423682196};
test_output[4220] = '{96.6512776079};
############ END DEBUG ############*/
test_input[33768:33775] = '{32'h4019dd98, 32'h419176f4, 32'h413d1a1f, 32'hc1f4638f, 32'hc1eca36a, 32'h42693f57, 32'hc26e74fb, 32'h41977ef2};
test_label[4221] = '{32'h419176f4};
test_output[4221] = '{32'h422083dd};
/*############ DEBUG ############
test_input[33768:33775] = '{2.40415004895, 18.1830833584, 11.8188772973, -30.5486129798, -29.5797916129, 58.3118548738, -59.6142370099, 18.9369852314};
test_label[4221] = '{18.1830833584};
test_output[4221] = '{40.1287715154};
############ END DEBUG ############*/
test_input[33776:33783] = '{32'hc25b2db9, 32'h42133de6, 32'h4251f026, 32'hc1f1ba1f, 32'hc23f75ea, 32'hc26819f3, 32'hc1489124, 32'hbf9aac0f};
test_label[4222] = '{32'hc23f75ea};
test_output[4222] = '{32'h42c8b308};
/*############ DEBUG ############
test_input[33776:33783] = '{-54.7946514315, 36.8104482676, 52.4845210931, -30.2158799391, -47.8651514954, -58.0253428488, -12.5354348704, -1.20837577664};
test_label[4222] = '{-47.8651514954};
test_output[4222] = '{100.349672744};
############ END DEBUG ############*/
test_input[33784:33791] = '{32'hc1a351bb, 32'hc2b94504, 32'hc27379df, 32'hc284efd6, 32'h42c0bbe8, 32'hc237ab45, 32'h4263f4bd, 32'h42b8ef38};
test_label[4223] = '{32'hc237ab45};
test_output[4223] = '{32'h430e4de7};
/*############ DEBUG ############
test_input[33784:33791] = '{-20.414907511, -92.6347931113, -60.8690147904, -66.4684282883, 96.36700561, -45.9172556127, 56.9890018227, 92.4672261962};
test_label[4223] = '{-45.9172556127};
test_output[4223] = '{142.304305367};
############ END DEBUG ############*/
test_input[33792:33799] = '{32'h42c20e97, 32'hc20d60d4, 32'hbfd5ff1a, 32'hc2b90631, 32'hc14effac, 32'hc10b8c96, 32'hc030e4df, 32'h4012edf0};
test_label[4224] = '{32'hc14effac};
test_output[4224] = '{32'h42dbee8d};
/*############ DEBUG ############
test_input[33792:33799] = '{97.0284989875, -35.3445605949, -1.67184762415, -92.512091002, -12.937420334, -8.72182253453, -2.76396914635, 2.29577246106};
test_label[4224] = '{-12.937420334};
test_output[4224] = '{109.965919322};
############ END DEBUG ############*/
test_input[33800:33807] = '{32'h428529b9, 32'hc29e9aa6, 32'h41e965fe, 32'hc26c855f, 32'h427e93ab, 32'h422eb40a, 32'h423b4be4, 32'h4217e1cd};
test_label[4225] = '{32'h427e93ab};
test_output[4225] = '{32'h403f4aa8};
/*############ DEBUG ############
test_input[33800:33807] = '{66.581487871, -79.3020451062, 29.1748000354, -59.1302462787, 63.6442086118, 43.6758181024, 46.8241138245, 37.9705066979};
test_label[4225] = '{63.6442086118};
test_output[4225] = '{2.98893176228};
############ END DEBUG ############*/
test_input[33808:33815] = '{32'hc2387b60, 32'h40fa165c, 32'hc17d042b, 32'h41a8700f, 32'h42a3242f, 32'h429ffd09, 32'h42ba423b, 32'h42530e89};
test_label[4226] = '{32'h42ba423b};
test_output[4226] = '{32'h374164fa};
/*############ DEBUG ############
test_input[33808:33815] = '{-46.1204852231, 7.81522948521, -15.8135172719, 21.0547153552, 81.5706686756, 79.9942096739, 93.1293575573, 52.7641944481};
test_label[4226] = '{93.1293575573};
test_output[4226] = '{1.15272066577e-05};
############ END DEBUG ############*/
test_input[33816:33823] = '{32'h425bdd5b, 32'hc136ae4b, 32'hc20b5118, 32'hc2a3bc80, 32'h42171637, 32'hc234c528, 32'hc194a239, 32'h4237e2d5};
test_label[4227] = '{32'h425bdd5b};
test_output[4227] = '{32'h3902205c};
/*############ DEBUG ############
test_input[33816:33823] = '{54.9661672336, -11.4175523489, -34.8291915477, -81.8681604262, 37.7716949428, -45.1925365672, -18.5792111161, 45.9715173389};
test_label[4227] = '{54.9661672336};
test_output[4227] = '{0.000124098211231};
############ END DEBUG ############*/
test_input[33824:33831] = '{32'h41dd5053, 32'hc1c7245e, 32'hc28937a0, 32'hc141d7cd, 32'h42078d6a, 32'h41af634a, 32'hc1370ff1, 32'h426849a2};
test_label[4228] = '{32'hc1c7245e};
test_output[4228] = '{32'h42a5ede8};
/*############ DEBUG ############
test_input[33824:33831] = '{27.6642204738, -24.8927579758, -68.6086437584, -12.1151855449, 33.8880992531, 21.923480212, -11.4413916199, 58.0719054413};
test_label[4228] = '{-24.8927579758};
test_output[4228] = '{82.9646634171};
############ END DEBUG ############*/
test_input[33832:33839] = '{32'h424b2040, 32'h428f6788, 32'h4145530d, 32'h42a08a4e, 32'hc204d291, 32'h4252b0ee, 32'hc22e9a10, 32'hc2adcded};
test_label[4229] = '{32'hc2adcded};
test_output[4229] = '{32'h43272c2a};
/*############ DEBUG ############
test_input[33832:33839] = '{50.7814953292, 71.7022073705, 12.3327758058, 80.2701238123, -33.2056321923, 52.6727841697, -43.6504528034, -86.9021960482};
test_label[4229] = '{-86.9021960482};
test_output[4229] = '{167.172509951};
############ END DEBUG ############*/
test_input[33840:33847] = '{32'h40a0fe0c, 32'hc2300cc4, 32'h4252ff18, 32'h4238076d, 32'h4040e67b, 32'hc1733e68, 32'h41c9eb8b, 32'hc20747f3};
test_label[4230] = '{32'h4238076d};
test_output[4230] = '{32'h40d7c703};
/*############ DEBUG ############
test_input[33840:33847] = '{5.03101169527, -44.0124646695, 52.7491166873, 46.007252871, 3.01406749028, -15.2027362842, 25.2400108776, -33.8202641507};
test_label[4230] = '{46.007252871};
test_output[4230] = '{6.74304356511};
############ END DEBUG ############*/
test_input[33848:33855] = '{32'hc254773b, 32'h415cbed3, 32'hc23eb8e6, 32'hc1babc1b, 32'h4201b9f5, 32'hc263d05c, 32'h4243640c, 32'h41d5e2de};
test_label[4231] = '{32'hc263d05c};
test_output[4231] = '{32'h42d39a34};
/*############ DEBUG ############
test_input[33848:33855] = '{-53.1164358514, 13.7965878786, -47.6805657058, -23.3418477694, 32.431598248, -56.9534748708, 48.8477009787, 26.7357748196};
test_label[4231] = '{-56.9534748708};
test_output[4231] = '{105.801175924};
############ END DEBUG ############*/
test_input[33856:33863] = '{32'hc25e32d7, 32'h3e8622f4, 32'h42a1307d, 32'h42462ef4, 32'hc113d2ac, 32'hc1a2c0b3, 32'hc2c167b3, 32'hc290ec39};
test_label[4232] = '{32'hc25e32d7};
test_output[4232] = '{32'h430824f4};
/*############ DEBUG ############
test_input[33856:33863] = '{-55.5496486513, 0.261985430825, 80.5947025054, 49.5458518188, -9.23893375791, -20.3440921948, -96.7025355949, -72.4613745699};
test_label[4232] = '{-55.5496486513};
test_output[4232] = '{136.144351157};
############ END DEBUG ############*/
test_input[33864:33871] = '{32'h42b8cd20, 32'hc11042a3, 32'hc2380529, 32'h421ae5f4, 32'hc10b8c44, 32'h42227978, 32'h4197260d, 32'h4230409e};
test_label[4233] = '{32'h4197260d};
test_output[4233] = '{32'h4293039c};
/*############ DEBUG ############
test_input[33864:33871] = '{92.4006310076, -9.01626829354, -46.0050383046, 38.7245639279, -8.72174419581, 40.6186203168, 18.8935786289, 44.0631026938};
test_label[4233] = '{18.8935786289};
test_output[4233] = '{73.5070523786};
############ END DEBUG ############*/
test_input[33872:33879] = '{32'h42b62ed3, 32'h40443d83, 32'hc2b00d45, 32'hc0bc72db, 32'hc220e6aa, 32'h42b9c348, 32'h42a126c5, 32'hc1845321};
test_label[4234] = '{32'h40443d83};
test_output[4234] = '{32'h42b3f06b};
/*############ DEBUG ############
test_input[33872:33879] = '{91.0914503527, 3.06625429545, -88.0259159702, -5.88902029026, -40.2252585199, 92.8814113736, 80.5757252053, -16.5405901742};
test_label[4234] = '{3.06625429545};
test_output[4234] = '{89.9695687557};
############ END DEBUG ############*/
test_input[33880:33887] = '{32'hc28a5d01, 32'hc0ccb7c9, 32'h40ab7b98, 32'h428fd8da, 32'h42922d41, 32'h41db1e9e, 32'h4284a474, 32'hc2823012};
test_label[4235] = '{32'h41db1e9e};
test_output[4235] = '{32'h4237e225};
/*############ DEBUG ############
test_input[33880:33887] = '{-69.1816501536, -6.39743492925, 5.35883696403, 71.9235381571, 73.0883848198, 27.3899494347, 66.3212012779, -65.0938858763};
test_label[4235] = '{27.3899494347};
test_output[4235] = '{45.9708424565};
############ END DEBUG ############*/
test_input[33888:33895] = '{32'hc2b6e6fa, 32'h4164f313, 32'hc2c5b04c, 32'hc211bdbe, 32'hc1b1148f, 32'h42244102, 32'h422b02a9, 32'h429c939f};
test_label[4236] = '{32'hc211bdbe};
test_output[4236] = '{32'h42e5727e};
/*############ DEBUG ############
test_input[33888:33895] = '{-91.4511284251, 14.309344367, -98.844331291, -36.4352948182, -22.1350391004, 41.0634837621, 42.7525987278, 78.2883196778};
test_label[4236] = '{-36.4352948182};
test_output[4236] = '{114.723614496};
############ END DEBUG ############*/
test_input[33896:33903] = '{32'h429bcf59, 32'h42b0e4fc, 32'h414b8d5c, 32'hc12f8d46, 32'h4036b0da, 32'hc2b523ef, 32'h428ca560, 32'hc2be2e4c};
test_label[4237] = '{32'h414b8d5c};
test_output[4237] = '{32'h42977354};
/*############ DEBUG ############
test_input[33896:33903] = '{77.9049741642, 88.4472353756, 12.7220116657, -10.9719904765, 2.85454415594, -90.5701808405, 70.3229992534, -95.0904233906};
test_label[4237] = '{12.7220116657};
test_output[4237] = '{75.7252501199};
############ END DEBUG ############*/
test_input[33904:33911] = '{32'h41317000, 32'hc28eb71e, 32'h41256f8a, 32'hc29df7bb, 32'h41fe0ce2, 32'hc25de5a9, 32'h4190916a, 32'hc284456e};
test_label[4238] = '{32'hc284456e};
test_output[4238] = '{32'h42c3c8a7};
/*############ DEBUG ############
test_input[33904:33911] = '{11.0898437237, -71.3576492644, 10.3397314503, -78.983845644, 31.7562909967, -55.474278317, 18.0710036181, -66.1356073322};
test_label[4238] = '{-66.1356073322};
test_output[4238] = '{97.8918994696};
############ END DEBUG ############*/
test_input[33912:33919] = '{32'hc10f97fe, 32'hc213457a, 32'h42884b0f, 32'h41cce565, 32'hc21b9050, 32'hc2917096, 32'hc1ac557e, 32'hc1454df5};
test_label[4239] = '{32'hc213457a};
test_output[4239] = '{32'h42d1edcc};
/*############ DEBUG ############
test_input[33912:33919] = '{-8.97460728911, -36.8178490158, 68.1466016302, 25.6120097933, -38.8909294866, -72.719895619, -21.5417433089, -12.331532403};
test_label[4239] = '{-36.8178490158};
test_output[4239] = '{104.964450646};
############ END DEBUG ############*/
test_input[33920:33927] = '{32'h422e6dd0, 32'h42c3446c, 32'h40f35c58, 32'hc2c63883, 32'h4277de80, 32'h42bab420, 32'h4206df4c, 32'h4123ac82};
test_label[4240] = '{32'hc2c63883};
test_output[4240] = '{32'h4344c1fb};
/*############ DEBUG ############
test_input[33920:33927] = '{43.6072391933, 97.6336371391, 7.60502247748, -99.1103767418, 61.9672852002, 93.3518036618, 33.7180625602, 10.2296159503};
test_label[4240] = '{-99.1103767418};
test_output[4240] = '{196.757736597};
############ END DEBUG ############*/
test_input[33928:33935] = '{32'hc2c23747, 32'h410814b7, 32'hc2840da6, 32'hc1116f12, 32'h408b0853, 32'hc2ac2e0f, 32'hc1a7a62c, 32'hc00ddbce};
test_label[4241] = '{32'hc2840da6};
test_output[4241] = '{32'h4295182d};
/*############ DEBUG ############
test_input[33928:33935] = '{-97.1079617688, 8.50505709814, -66.0266553231, -9.08961711856, 4.34476629341, -86.0899591965, -20.9561395084, -2.21654078178};
test_label[4241] = '{-66.0266553231};
test_output[4241] = '{74.5472167121};
############ END DEBUG ############*/
test_input[33936:33943] = '{32'hc2a1c6bf, 32'h4065f9e7, 32'hc23a3edb, 32'h42908d72, 32'hc2023355, 32'h422ad3cd, 32'h4287b940, 32'h4285743b};
test_label[4242] = '{32'h422ad3cd};
test_output[4242] = '{32'h41ecaeae};
/*############ DEBUG ############
test_input[33936:33943] = '{-80.8881759529, 3.59337773354, -46.5613836979, 72.2762623926, -32.5501275895, 42.7068353149, 67.8618133638, 66.7270116848};
test_label[4242] = '{42.7068353149};
test_output[4242] = '{29.5852921502};
############ END DEBUG ############*/
test_input[33944:33951] = '{32'hc1e36fcf, 32'hc13d612f, 32'h428e3896, 32'h4019966e, 32'h410b2b84, 32'hc28b7b3d, 32'hc29a5baa, 32'hc1916353};
test_label[4243] = '{32'hc28b7b3d};
test_output[4243] = '{32'h430cd9e9};
/*############ DEBUG ############
test_input[33944:33951] = '{-28.4295937446, -11.8362268469, 71.1105196871, 2.39980640957, 8.69812348795, -69.7406972225, -77.1790338311, -18.1734977553};
test_label[4243] = '{-69.7406972225};
test_output[4243] = '{140.85121691};
############ END DEBUG ############*/
test_input[33952:33959] = '{32'h42b745cc, 32'h413e83fe, 32'hc2321e24, 32'h420596f1, 32'h42ba97d6, 32'hc12517f5, 32'hc28ea6be, 32'h4189f0fb};
test_label[4244] = '{32'h413e83fe};
test_output[4244] = '{32'h42a32071};
/*############ DEBUG ############
test_input[33952:33959] = '{91.6363198197, 11.9072250574, -44.5294350103, 33.3974035952, 93.2965529335, -10.3183484131, -71.3256721005, 17.2426666376};
test_label[4244] = '{11.9072250574};
test_output[4244] = '{81.5633607274};
############ END DEBUG ############*/
test_input[33960:33967] = '{32'hc2a04e79, 32'h425fe511, 32'hc1f640b5, 32'h42688f8b, 32'hc239a9bf, 32'h42a80f97, 32'hc1c6510a, 32'hc2917a20};
test_label[4245] = '{32'hc239a9bf};
test_output[4245] = '{32'h4302723b};
/*############ DEBUG ############
test_input[33960:33967] = '{-80.1532676102, 55.9736962487, -30.781596082, 58.1401804788, -46.4157675184, 84.0304503362, -24.7895706648, -72.7385218622};
test_label[4245] = '{-46.4157675184};
test_output[4245] = '{130.446217855};
############ END DEBUG ############*/
test_input[33968:33975] = '{32'h42031f82, 32'h42b99b6a, 32'h42af5443, 32'h42a95a25, 32'hc2bc74cb, 32'hc2555a9d, 32'h412649f1, 32'hc2a28236};
test_label[4246] = '{32'h42a95a25};
test_output[4246] = '{32'h4102234a};
/*############ DEBUG ############
test_input[33968:33975] = '{32.7807695174, 92.8035413752, 87.6645720206, 84.6760663774, -94.2281139874, -53.3384893753, 10.3930519352, -81.2543188365};
test_label[4246] = '{84.6760663774};
test_output[4246] = '{8.13361515136};
############ END DEBUG ############*/
test_input[33976:33983] = '{32'h42b77209, 32'hc2c4f1e9, 32'hc1240b11, 32'hc16469e5, 32'hc2bc8800, 32'h41e6794f, 32'h42a6702e, 32'h4174b1d6};
test_label[4247] = '{32'h42a6702e};
test_output[4247] = '{32'h41080fa9};
/*############ DEBUG ############
test_input[33976:33983] = '{91.7227226834, -98.4724828634, -10.2527015592, -14.2758532691, -94.2656237923, 28.8092318868, 83.2191021183, 15.2934167889};
test_label[4247] = '{83.2191021183};
test_output[4247] = '{8.50382327766};
############ END DEBUG ############*/
test_input[33984:33991] = '{32'h429666a4, 32'hc15bd9cc, 32'h402152f7, 32'h41c1787e, 32'h426e648b, 32'h41b590a7, 32'h42418c57, 32'hc29cddcc};
test_label[4248] = '{32'h429666a4};
test_output[4248] = '{32'h3433dabf};
/*############ DEBUG ############
test_input[33984:33991] = '{75.2004688712, -13.7406734219, 2.52068874424, 24.1838345543, 59.5981881129, 22.6956302167, 48.3870504601, -78.433196248};
test_label[4248] = '{75.2004688712};
test_output[4248] = '{1.67502540433e-07};
############ END DEBUG ############*/
test_input[33992:33999] = '{32'h42c25967, 32'h42a1c1d7, 32'hc238ac78, 32'h4124d1ec, 32'hc29103eb, 32'hc2c503f6, 32'hc1866811, 32'hc23fac8e};
test_label[4249] = '{32'h42a1c1d7};
test_output[4249] = '{32'h41825e3f};
/*############ DEBUG ############
test_input[33992:33999] = '{97.1746141466, 80.8785959794, -46.1684278451, 10.3012508085, -72.5076487186, -98.5077380885, -16.8008142742, -47.9185118719};
test_label[4249] = '{80.8785959794};
test_output[4249] = '{16.2960182509};
############ END DEBUG ############*/
test_input[34000:34007] = '{32'h419a9622, 32'hc1d245cc, 32'hc0aa4125, 32'hc2a9bfea, 32'h42ad738a, 32'hc2834cb1, 32'h417d0cc1, 32'h41f088f7};
test_label[4250] = '{32'h419a9622};
test_output[4250] = '{32'h4286ce01};
/*############ DEBUG ############
test_input[34000:34007] = '{19.32330637, -26.2840802872, -5.32045212067, -84.8748349566, 86.7256593146, -65.6497916771, 15.8156133283, 30.0668774466};
test_label[4250] = '{19.32330637};
test_output[4250] = '{67.4023529446};
############ END DEBUG ############*/
test_input[34008:34015] = '{32'hc1329026, 32'h42388e9c, 32'h4036dd8f, 32'h4219e58d, 32'hc18bfc1c, 32'h41a2aae8, 32'h429f6e54, 32'hc2c79dbc};
test_label[4251] = '{32'h4036dd8f};
test_output[4251] = '{32'h4299b768};
/*############ DEBUG ############
test_input[34008:34015] = '{-11.1601924075, 46.1392664984, 2.85727295774, 38.4741716659, -17.4981010355, 20.3334494002, 79.715488358, -99.8080724859};
test_label[4251] = '{2.85727295774};
test_output[4251] = '{76.8582154003};
############ END DEBUG ############*/
test_input[34016:34023] = '{32'h41a15420, 32'h42accccc, 32'hc286bfb0, 32'h42b938e5, 32'h41cfb247, 32'h42365122, 32'hc142f9c0, 32'hc29b7c31};
test_label[4252] = '{32'h41cfb247};
test_output[4252] = '{32'h42854d5a};
/*############ DEBUG ############
test_input[34016:34023] = '{20.1660770592, 86.399995203, -67.3743893703, 92.6111185888, 25.9620499195, 45.5792309148, -12.1859744502, -77.7425606658};
test_label[4252] = '{25.9620499195};
test_output[4252] = '{66.6510736396};
############ END DEBUG ############*/
test_input[34024:34031] = '{32'hc2a25b0a, 32'hc1ab90e0, 32'hc150e905, 32'hc0989e9b, 32'hc271bed9, 32'h42bef88f, 32'h42067da4, 32'hc20c139e};
test_label[4253] = '{32'hc20c139e};
test_output[4253] = '{32'h4302812f};
/*############ DEBUG ############
test_input[34024:34031] = '{-81.1778083036, -21.4457392606, -13.0568894805, -4.76936108007, -60.436375088, 95.4854694065, 33.622695511, -35.0191583229};
test_label[4253] = '{-35.0191583229};
test_output[4253] = '{130.504627729};
############ END DEBUG ############*/
test_input[34032:34039] = '{32'hc20d9a81, 32'h41f071d2, 32'h42a4a2ca, 32'hc28a461b, 32'hc25cea1d, 32'hbffb6b6b, 32'h414eae50, 32'hc16fb8b4};
test_label[4254] = '{32'h42a4a2ca};
test_output[4254] = '{32'h80000000};
/*############ DEBUG ############
test_input[34032:34039] = '{-35.4008839276, 30.0555758489, 82.3179504116, -69.1369271741, -55.2286246278, -1.96421567718, 12.9175568823, -14.9825930608};
test_label[4254] = '{82.3179504116};
test_output[4254] = '{-0.0};
############ END DEBUG ############*/
test_input[34040:34047] = '{32'h4285fcd5, 32'hc1e55e02, 32'h414a3636, 32'h418f4083, 32'h420680ba, 32'hc2868866, 32'h42a609f3, 32'h42925371};
test_label[4255] = '{32'h414a3636};
test_output[4255] = '{32'h428cc333};
/*############ DEBUG ############
test_input[34040:34047] = '{66.9938150287, -28.6709029349, 12.6382350388, 17.9065000663, 33.6257092505, -67.2664040606, 83.0194332539, 73.1629750798};
test_label[4255] = '{12.6382350388};
test_output[4255] = '{70.381250731};
############ END DEBUG ############*/
test_input[34048:34055] = '{32'hc2c29040, 32'h429ed434, 32'h427a5960, 32'h4272ecac, 32'h4217486e, 32'hc2516802, 32'hc18d1b08, 32'h425df25d};
test_label[4256] = '{32'h429ed434};
test_output[4256] = '{32'h33748e77};
/*############ DEBUG ############
test_input[34048:34055] = '{-97.2817383367, 79.4144583929, 62.5872811612, 60.7311233655, 37.8207314924, -52.3515711009, -17.6381987099, 55.4866834268};
test_label[4256] = '{79.4144583929};
test_output[4256] = '{5.6940248361e-08};
############ END DEBUG ############*/
test_input[34056:34063] = '{32'h423a76e7, 32'hc1fb4e81, 32'h42ad5794, 32'hc0d595de, 32'h41e930ea, 32'hc2bc3ba4, 32'h426a17aa, 32'h42025412};
test_label[4257] = '{32'h423a76e7};
test_output[4257] = '{32'h42203842};
/*############ DEBUG ############
test_input[34056:34063] = '{46.616113852, -31.4133319231, 86.6710530701, -6.67454447375, 29.1488835358, -94.1164841281, 58.5231110595, 32.5820987753};
test_label[4257] = '{46.616113852};
test_output[4257] = '{40.0549392181};
############ END DEBUG ############*/
test_input[34064:34071] = '{32'hc1e57748, 32'hc245d80e, 32'h429e6210, 32'h42b7fa33, 32'hc237d599, 32'h42b4cb0d, 32'h424296e5, 32'hc0807656};
test_label[4258] = '{32'hc1e57748};
test_output[4258] = '{32'h42f1b6dd};
/*############ DEBUG ############
test_input[34064:34071] = '{-28.6832423282, -49.4609921383, 79.1915306877, 91.9886735589, -45.9585912691, 90.3965801075, 48.6473563721, -4.01444530835};
test_label[4258] = '{-28.6832423282};
test_output[4258] = '{120.85715146};
############ END DEBUG ############*/
test_input[34072:34079] = '{32'hc2bb385e, 32'h422d9c1b, 32'h42bf3982, 32'hc29c1804, 32'hc215d92f, 32'hc0bced40, 32'h41e8df68, 32'hc01d59b6};
test_label[4259] = '{32'hc215d92f};
test_output[4259] = '{32'h4305130d};
/*############ DEBUG ############
test_input[34072:34079] = '{-93.6100897603, 43.4024452412, 95.6123203348, -78.046905065, -37.4620945105, -5.9039610384, 29.1090857741, -2.45860042687};
test_label[4259] = '{-37.4620945105};
test_output[4259] = '{133.074414845};
############ END DEBUG ############*/
test_input[34080:34087] = '{32'hc20cf9a3, 32'hc1f51da3, 32'hc1a97957, 32'hc2bf8bef, 32'h4241e969, 32'hc1db926a, 32'h42407346, 32'h42bf4162};
test_label[4260] = '{32'h42bf4162};
test_output[4260] = '{32'h80000000};
/*############ DEBUG ############
test_input[34080:34087] = '{-35.2437873788, -30.6394709623, -21.1842488464, -95.7733059437, 48.4779389266, -27.4464912638, 48.1125710775, 95.6276995959};
test_label[4260] = '{95.6276995959};
test_output[4260] = '{-0.0};
############ END DEBUG ############*/
test_input[34088:34095] = '{32'hc2abe750, 32'h42878c12, 32'hc2bec59c, 32'hc16a8c3b, 32'hc298ccf3, 32'hc2c5a4db, 32'hc2711745, 32'hc1093cf2};
test_label[4261] = '{32'hc2711745};
test_output[4261] = '{32'h43000bda};
/*############ DEBUG ############
test_input[34088:34095] = '{-85.9517836325, 67.77357336, -95.3859561073, -14.6592358598, -76.4002898308, -98.821982332, -60.2727246423, -8.57737953356};
test_label[4261] = '{-60.2727246423};
test_output[4261] = '{128.046298002};
############ END DEBUG ############*/
test_input[34096:34103] = '{32'hc285cfd3, 32'hc19c34ef, 32'h41863eb6, 32'h419d1960, 32'h429699b1, 32'hc1b65300, 32'hc287e1e7, 32'h4195d87b};
test_label[4262] = '{32'hc19c34ef};
test_output[4262] = '{32'h42bda6ec};
/*############ DEBUG ############
test_input[34096:34103] = '{-66.9059087038, -19.5258470002, 16.780620799, 19.6373906031, 75.3001757025, -22.7905269809, -67.9412123265, 18.7307025153};
test_label[4262] = '{-19.5258470002};
test_output[4262] = '{94.8260227027};
############ END DEBUG ############*/
test_input[34104:34111] = '{32'h42c13cf6, 32'hc2346398, 32'hc246b14c, 32'hc2b6421b, 32'h419309db, 32'hc24790fb, 32'h42bd21ef, 32'hc2718a09};
test_label[4263] = '{32'h419309db};
test_output[4263] = '{32'h429cb856};
/*############ DEBUG ############
test_input[34104:34111] = '{96.6190633114, -45.0972589134, -49.6731408943, -91.1291132893, 18.3798125006, -49.8915822541, 94.5662737958, -60.384801238};
test_label[4263] = '{18.3798125006};
test_output[4263] = '{78.3600305039};
############ END DEBUG ############*/
test_input[34112:34119] = '{32'h42987570, 32'hc1b7e4ea, 32'h42ba4450, 32'h42c12bb4, 32'h4053e5c3, 32'hc292a250, 32'h4204b8cc, 32'hc2b6c409};
test_label[4264] = '{32'hc292a250};
test_output[4264] = '{32'h4329eefe};
/*############ DEBUG ############
test_input[34112:34119] = '{76.2293679919, -22.9867742605, 93.1334210427, 96.5853545874, 3.31089856389, -73.3170142381, 33.1804658523, -91.3828830126};
test_label[4264] = '{-73.3170142381};
test_output[4264] = '{169.93356155};
############ END DEBUG ############*/
test_input[34120:34127] = '{32'hc1c4cffe, 32'h42983653, 32'h425301c0, 32'h42b195a0, 32'hc2842759, 32'h42973911, 32'hc2c470b8, 32'hc1c52ff9};
test_label[4265] = '{32'h42983653};
test_output[4265] = '{32'h414afa6a};
/*############ DEBUG ############
test_input[34120:34127] = '{-24.601558517, 76.106103455, 52.7517097705, 88.7922349395, -66.0768473401, 75.6114570876, -98.2201550758, -24.6484247196};
test_label[4265] = '{76.106103455};
test_output[4265] = '{12.6861364647};
############ END DEBUG ############*/
test_input[34128:34135] = '{32'hc2bd7c88, 32'h4200c463, 32'hc2007e8e, 32'h42a43edd, 32'h421ea11d, 32'hbff8eff6, 32'hc25b4ad5, 32'h42bab9b7};
test_label[4266] = '{32'hc25b4ad5};
test_output[4266] = '{32'h43142f91};
/*############ DEBUG ############
test_input[34128:34135] = '{-94.7432245153, 32.1917850245, -32.1235890531, 82.1227783179, 39.6573364061, -1.94482299049, -54.8230762537, 93.3627237429};
test_label[4266] = '{-54.8230762537};
test_output[4266] = '{148.185813135};
############ END DEBUG ############*/
test_input[34136:34143] = '{32'h42a37fda, 32'h42c1eccf, 32'h4210c1be, 32'h429c463b, 32'hc285a5e5, 32'h42a992b1, 32'hc22bc12e, 32'hc15ad5f6};
test_label[4267] = '{32'h42a992b1};
test_output[4267] = '{32'h4142d0fa};
/*############ DEBUG ############
test_input[34136:34143] = '{81.7497072193, 96.9625188932, 36.1892023446, 78.1371674629, -66.8240133617, 84.7865048976, -42.9386530334, -13.6772364099};
test_label[4267] = '{84.7865048976};
test_output[4267] = '{12.1760194021};
############ END DEBUG ############*/
test_input[34144:34151] = '{32'h41cc1128, 32'hc2c4d5e9, 32'h42b1b80c, 32'hc2add866, 32'hc2a965a1, 32'h42bd0b25, 32'h422bfaa9, 32'hc27c56ae};
test_label[4268] = '{32'hc2add866};
test_output[4268] = '{32'h433572a9};
/*############ DEBUG ############
test_input[34144:34151] = '{25.5083767475, -98.4177896976, 88.8594632808, -86.9226531117, -84.6984971008, 94.5217632794, 42.9947861624, -63.084649455};
test_label[4268] = '{-86.9226531117};
test_output[4268] = '{181.447884885};
############ END DEBUG ############*/
test_input[34152:34159] = '{32'hc231231b, 32'hc1480746, 32'h421b1f07, 32'h42b48c8a, 32'hc2a94f9d, 32'hc2a0978d, 32'h42b4773e, 32'hc23e022b};
test_label[4269] = '{32'hc2a94f9d};
test_output[4269] = '{32'h432f9a41};
/*############ DEBUG ############
test_input[34152:34159] = '{-44.2842830315, -12.5017755333, 38.7802986352, 90.2744869705, -84.6554925348, -80.2959994408, 90.232896575, -47.5021164459};
test_label[4269] = '{-84.6554925348};
test_output[4269] = '{175.602547693};
############ END DEBUG ############*/
test_input[34160:34167] = '{32'h420ef731, 32'hc1e8b212, 32'hc124a165, 32'h408cc3a1, 32'h427744c3, 32'hc2801897, 32'h421a7a64, 32'hc2a8c505};
test_label[4270] = '{32'hc2801897};
test_output[4270] = '{32'h42fbbaf8};
/*############ DEBUG ############
test_input[34160:34167] = '{35.7413959584, -29.0869475067, -10.2894027506, 4.39888048764, 61.8171511041, -64.0480239436, 38.6195204043, -84.3848003161};
test_label[4270] = '{-64.0480239436};
test_output[4270] = '{125.865175048};
############ END DEBUG ############*/
test_input[34168:34175] = '{32'hc2b9efde, 32'h4226f981, 32'hc29e70be, 32'hc2a4a6d5, 32'hc2c6e73e, 32'hc26c4aff, 32'h424c2e15, 32'h4223ba24};
test_label[4271] = '{32'h4226f981};
test_output[4271] = '{32'h4114d2d8};
/*############ DEBUG ############
test_input[34168:34175] = '{-92.9684909652, 41.7436577184, -79.220198415, -82.3258404101, -99.4516424921, -59.0732365107, 51.0450012948, 40.9317760888};
test_label[4271] = '{41.7436577184};
test_output[4271] = '{9.30147540903};
############ END DEBUG ############*/
test_input[34176:34183] = '{32'hc202333f, 32'h4119b826, 32'hbc957b9f, 32'h42a00e9e, 32'hc28e08a2, 32'h40e85451, 32'h42180255, 32'h409a1169};
test_label[4272] = '{32'h42180255};
test_output[4272] = '{32'h42281ae8};
/*############ DEBUG ############
test_input[34176:34183] = '{-32.5500433581, 9.60745784975, -0.0182474242405, 80.0285502849, -71.0168616773, 7.26029242967, 38.0022761916, 4.81462545506};
test_label[4272] = '{38.0022761916};
test_output[4272] = '{42.0262740933};
############ END DEBUG ############*/
test_input[34184:34191] = '{32'hbec5eb70, 32'hbd97e587, 32'h42c13ef5, 32'hc2bf1707, 32'h42c515b8, 32'h42b50cea, 32'hc2af1cf6, 32'hc24be408};
test_label[4273] = '{32'hbd97e587};
test_output[4273] = '{32'h42c581eb};
/*############ DEBUG ############
test_input[34184:34191] = '{-0.386561882778, -0.0741682588418, 96.6229600659, -95.5449790159, 98.5424167255, 90.5252197315, -87.5565629128, -50.972686051};
test_label[4273] = '{-0.0741682588418};
test_output[4273] = '{98.7537491069};
############ END DEBUG ############*/
test_input[34192:34199] = '{32'h42553739, 32'hc22f447c, 32'h41208bb8, 32'h416bf20e, 32'hc2364226, 32'h42bd6fda, 32'hc288abcf, 32'hc29eae4a};
test_label[4274] = '{32'h42bd6fda};
test_output[4274] = '{32'h80000000};
/*############ DEBUG ############
test_input[34192:34199] = '{53.3039292606, -43.8168785733, 10.0341109896, 14.7465952527, -45.5645991111, 94.7184602068, -68.3355621227, -79.3404053333};
test_label[4274] = '{94.7184602068};
test_output[4274] = '{-0.0};
############ END DEBUG ############*/
test_input[34200:34207] = '{32'h41fa7014, 32'hc2a7279b, 32'hc23147a5, 32'h428a1b1e, 32'hc287a043, 32'h41d3aa98, 32'h42938f34, 32'h42a22fd7};
test_label[4275] = '{32'h41d3aa98};
test_output[4275] = '{32'h425a8b11};
/*############ DEBUG ############
test_input[34200:34207] = '{31.3047262281, -83.5773546137, -44.3199646879, 69.0529605957, -67.8130114564, 26.4582980781, 73.7796934581, 81.0934344432};
test_label[4275] = '{26.4582980781};
test_output[4275] = '{54.6358083595};
############ END DEBUG ############*/
test_input[34208:34215] = '{32'hc205870f, 32'h42863c24, 32'hc2146d3e, 32'h3f0d27b8, 32'hc2785037, 32'hc20cf5ce, 32'hc2160501, 32'h4295cc38};
test_label[4276] = '{32'hc2785037};
test_output[4276] = '{32'h4308fa45};
/*############ DEBUG ############
test_input[34208:34215] = '{-33.3818930271, 67.1174585746, -37.1066832304, 0.551387292033, -62.078334847, -35.2400443336, -37.5048863612, 74.8988640838};
test_label[4276] = '{-62.078334847};
test_output[4276] = '{136.977616269};
############ END DEBUG ############*/
test_input[34216:34223] = '{32'hc239b055, 32'hc28d979c, 32'h429f8139, 32'h415196bf, 32'h42b1d206, 32'hc26391b0, 32'hc1aa28cd, 32'h41b6c634};
test_label[4277] = '{32'hc239b055};
test_output[4277] = '{32'h4307551f};
/*############ DEBUG ############
test_input[34216:34223] = '{-46.4221999074, -70.7961114943, 79.7523888908, 13.0993032013, 88.9101990164, -56.892273528, -21.2699222204, 22.8467784398};
test_label[4277] = '{-46.4221999074};
test_output[4277] = '{135.332504312};
############ END DEBUG ############*/
test_input[34224:34231] = '{32'hc28a0eac, 32'h411270e8, 32'h41f5d4ad, 32'hc1330376, 32'h41ba6472, 32'h40b3793b, 32'hc25cae92, 32'hc1cd0086};
test_label[4278] = '{32'h41f5d4ad};
test_output[4278] = '{32'h3a1b7c58};
/*############ DEBUG ############
test_input[34224:34231] = '{-69.0286552694, 9.15256461176, 30.728845804, -11.188344813, 23.2990462337, 5.60854887674, -55.1704806047, -25.6252551781};
test_label[4278] = '{30.728845804};
test_output[4278] = '{0.000593130917726};
############ END DEBUG ############*/
test_input[34232:34239] = '{32'h421d22a9, 32'hc114afca, 32'hc2978289, 32'hc28863f7, 32'hc28dc478, 32'h4240c4ed, 32'h429b265a, 32'hc0862c5a};
test_label[4279] = '{32'hc0862c5a};
test_output[4279] = '{32'h42a38920};
/*############ DEBUG ############
test_input[34232:34239] = '{39.2838467348, -9.29291724022, -75.7549534445, -68.1952468481, -70.8837254576, 48.192309099, 77.5749044816, -4.19291408388};
test_label[4279] = '{-4.19291408388};
test_output[4279] = '{81.7678185655};
############ END DEBUG ############*/
test_input[34240:34247] = '{32'hc28605cb, 32'h419618c0, 32'hc226506a, 32'h42c37f84, 32'h42c4377f, 32'h41072cd3, 32'hc28872c7, 32'h419c87e7};
test_label[4280] = '{32'hc226506a};
test_output[4280] = '{32'h430c376a};
/*############ DEBUG ############
test_input[34240:34247] = '{-67.0113159683, 18.7620855225, -41.5785295525, 97.7490577527, 98.1083922108, 8.44844348516, -68.2241713746, 19.566358733};
test_label[4280] = '{-41.5785295525};
test_output[4280] = '{140.216455777};
############ END DEBUG ############*/
test_input[34248:34255] = '{32'h41713e08, 32'h425da804, 32'hc2940d26, 32'hc2263674, 32'h42bd7cd7, 32'hc2b04b73, 32'hc2265643, 32'hc291d174};
test_label[4281] = '{32'h425da804};
test_output[4281] = '{32'h421d51aa};
/*############ DEBUG ############
test_input[34248:34255] = '{15.0776443785, 55.4140769203, -74.0256830636, -41.5531784195, 94.7438268963, -88.1473645501, -41.5842395486, -72.9090901068};
test_label[4281] = '{55.4140769203};
test_output[4281] = '{39.329749976};
############ END DEBUG ############*/
test_input[34256:34263] = '{32'h420ba1d3, 32'h4285ca80, 32'hc19b9fe5, 32'hc2308552, 32'hc2085981, 32'h4280ee29, 32'h420e37d1, 32'hc21d5a5e};
test_label[4282] = '{32'hc2308552};
test_output[4282] = '{32'h42de3859};
/*############ DEBUG ############
test_input[34256:34263] = '{34.9080302594, 66.8955095991, -19.4530732929, -44.1301974922, -34.0874047085, 64.4651531006, 35.554509023, -39.338249525};
test_label[4282] = '{-44.1301974922};
test_output[4282] = '{111.110053252};
############ END DEBUG ############*/
test_input[34264:34271] = '{32'hc1ea236e, 32'h42be3be9, 32'hc1f85954, 32'h414ae36d, 32'h42b226ed, 32'h4285aa37, 32'h427851d6, 32'hc1ae4c0d};
test_label[4283] = '{32'h414ae36d};
test_output[4283] = '{32'h42a4e0b3};
/*############ DEBUG ############
test_input[34264:34271] = '{-29.2673001315, 95.1170125732, -31.0436180875, 12.6805234607, 89.0760262284, 66.8324493254, 62.0799172148, -21.7871332834};
test_label[4283] = '{12.6805234607};
test_output[4283] = '{82.4388654978};
############ END DEBUG ############*/
test_input[34272:34279] = '{32'h405bc201, 32'hc0eece54, 32'hc2209d1a, 32'hc293cfd7, 32'hc29f85e1, 32'h429f9d28, 32'hc23ea44b, 32'hc2af2e2c};
test_label[4284] = '{32'hc0eece54};
test_output[4284] = '{32'h42ae8a0d};
/*############ DEBUG ############
test_input[34272:34279] = '{3.43371607325, -7.46268668301, -40.1534204374, -73.9059387823, -79.7614795335, 79.806946635, -47.6604434472, -87.5901764391};
test_label[4284] = '{-7.46268668301};
test_output[4284] = '{87.269633318};
############ END DEBUG ############*/
test_input[34280:34287] = '{32'h42b41d15, 32'h428c6279, 32'h42847a79, 32'h42950549, 32'h422e64a9, 32'h42aaa1d9, 32'hc0307e94, 32'hc2b4c88b};
test_label[4285] = '{32'h428c6279};
test_output[4285] = '{32'h419efc3d};
/*############ DEBUG ############
test_input[34280:34287] = '{90.0567998741, 70.1923316653, 66.2392010236, 74.5103197822, 43.5983022575, 85.3161092646, -2.75772566686, -90.3916880931};
test_label[4285] = '{70.1923316653};
test_output[4285] = '{19.8731630913};
############ END DEBUG ############*/
test_input[34288:34295] = '{32'hc1810b3c, 32'hc285eb36, 32'hc225e70a, 32'hc2afa946, 32'hc1394396, 32'hc0a9aad7, 32'hc18ab0db, 32'h42b990ab};
test_label[4286] = '{32'hc0a9aad7};
test_output[4286] = '{32'h42c42b58};
/*############ DEBUG ############
test_input[34288:34295] = '{-16.1304864749, -66.9593996353, -41.4756226031, -87.8306106206, -11.5790002143, -5.30210437434, -17.3363558258, 92.7825534965};
test_label[4286] = '{-5.30210437434};
test_output[4286] = '{98.0846578708};
############ END DEBUG ############*/
test_input[34296:34303] = '{32'hc11ddea3, 32'hc1e52be7, 32'h423e6ec9, 32'hc22f841b, 32'hc1cb9378, 32'hc2c7110b, 32'h42c7e4ab, 32'h42206bf8};
test_label[4287] = '{32'hc2c7110b};
test_output[4287] = '{32'h43477adb};
/*############ DEBUG ############
test_input[34296:34303] = '{-9.86685472212, -28.6464358751, 47.6081879197, -43.8790097227, -25.4470069442, -99.533285525, 99.9466183092, 40.1054389172};
test_label[4287] = '{-99.533285525};
test_output[4287] = '{199.479903834};
############ END DEBUG ############*/
test_input[34304:34311] = '{32'h429c7eac, 32'h41d4b651, 32'hc1c84e3b, 32'hc27b4619, 32'h42199692, 32'hc29d3174, 32'h4163118f, 32'hc22199ec};
test_label[4288] = '{32'hc29d3174};
test_output[4288] = '{32'h431cd810};
/*############ DEBUG ############
test_input[34304:34311] = '{78.2474068768, 26.5890212094, -25.0381977939, -62.8184554652, 38.3970414467, -78.5965894392, 14.1917869881, -40.4003148043};
test_label[4288] = '{-78.5965894392};
test_output[4288] = '{156.843996316};
############ END DEBUG ############*/
test_input[34312:34319] = '{32'h428a183d, 32'h42aacc0d, 32'hc21c520a, 32'hc28269c3, 32'hc1fc59c8, 32'h42a606be, 32'h426273ec, 32'h410dd870};
test_label[4289] = '{32'h42aacc0d};
test_output[4289] = '{32'h3db459ae};
/*############ DEBUG ############
test_input[34312:34319] = '{69.0473392544, 85.3985363796, -39.0801165745, -65.2065621249, -31.5438377245, 83.0131715877, 56.6132053302, 8.86534076668};
test_label[4289] = '{85.3985363796};
test_output[4289] = '{0.0880616742003};
############ END DEBUG ############*/
test_input[34320:34327] = '{32'hc1a9e50f, 32'hc2372343, 32'hc2ba2fa6, 32'hc1e64041, 32'h42271443, 32'h42b9fe3e, 32'hc0ec5bea, 32'h41ff68cf};
test_label[4290] = '{32'hc2ba2fa6};
test_output[4290] = '{32'h433a16f2};
/*############ DEBUG ############
test_input[34320:34327] = '{-21.2368459302, -45.7844358529, -93.0930619582, -28.7813746505, 41.7697878911, 92.9965648038, -7.38622006066, 31.9261752963};
test_label[4290] = '{-93.0930619582};
test_output[4290] = '{186.089626762};
############ END DEBUG ############*/
test_input[34328:34335] = '{32'hc2a9b9f5, 32'h4072308b, 32'h41e548c4, 32'h42a8e2d9, 32'h42a373a1, 32'hc28ab883, 32'hc10a3d2c, 32'h422a0af6};
test_label[4291] = '{32'h41e548c4};
test_output[4291] = '{32'h425f62d0};
/*############ DEBUG ############
test_input[34328:34335] = '{-84.8631983049, 3.78421280508, 28.6605298899, 84.4430597641, 81.7258377209, -69.3603718492, -8.63993472872, 42.5107045997};
test_label[4291] = '{28.6605298899};
test_output[4291] = '{55.8464976131};
############ END DEBUG ############*/
test_input[34336:34343] = '{32'hc28324e7, 32'hc2b48246, 32'hc25717a9, 32'hc013be19, 32'h41d9df47, 32'h424c9dc0, 32'hc2ac3fcb, 32'h42c19429};
test_label[4292] = '{32'hc013be19};
test_output[4292] = '{32'h42c6321a};
/*############ DEBUG ############
test_input[34336:34343] = '{-65.5720736232, -90.254437953, -53.7731044674, -2.3084776568, 27.2340219949, 51.154053397, -86.1245927646, 96.7893741704};
test_label[4292] = '{-2.3084776568};
test_output[4292] = '{99.0978518272};
############ END DEBUG ############*/
test_input[34344:34351] = '{32'h425bb50b, 32'hc25924b3, 32'hc2b42b14, 32'hc2330874, 32'h429c5d38, 32'h4210b919, 32'h42102088, 32'hc24c5635};
test_label[4293] = '{32'h429c5d38};
test_output[4293] = '{32'h2eaed260};
/*############ DEBUG ############
test_input[34344:34351] = '{54.9268006465, -54.2858378906, -90.0841382656, -44.7582554242, 78.1820685222, 36.1807588239, 36.0317689206, -51.0841877437};
test_label[4293] = '{78.1820685222};
test_output[4293] = '{7.94997401275e-11};
############ END DEBUG ############*/
test_input[34352:34359] = '{32'h42a5c6a0, 32'hc266e988, 32'h420f5c47, 32'h4290c846, 32'hc24926af, 32'h42a9a1f1, 32'h429e42db, 32'h42bee536};
test_label[4294] = '{32'hc24926af};
test_output[4294] = '{32'h4311bc48};
/*############ DEBUG ############
test_input[34352:34359] = '{82.8879375286, -57.728059297, 35.8401164664, 72.391160574, -50.2877757946, 84.8162933968, 79.1305753596, 95.4476739622};
test_label[4294] = '{-50.2877757946};
test_output[4294] = '{145.735477495};
############ END DEBUG ############*/
test_input[34360:34367] = '{32'h420674db, 32'h41ade7a7, 32'hc290af4f, 32'h421c9bee, 32'h41941b8d, 32'h424f91e2, 32'h42359e98, 32'h41ba54ee};
test_label[4295] = '{32'h41ba54ee};
test_output[4295] = '{32'h41e4d1f6};
/*############ DEBUG ############
test_input[34360:34367] = '{33.6141152486, 21.7381118129, -72.3423977528, 39.1522757244, 18.5134518806, 51.8924653215, 45.4048763625, 23.2914698047};
test_label[4295] = '{23.2914698047};
test_output[4295] = '{28.602519512};
############ END DEBUG ############*/
test_input[34368:34375] = '{32'hc28e62af, 32'h42902dcb, 32'h42078b92, 32'hc25960bd, 32'hc27d2be4, 32'h42c7917e, 32'h41064976, 32'h42168ea7};
test_label[4296] = '{32'hc28e62af};
test_output[4296] = '{32'h432afa16};
/*############ DEBUG ############
test_input[34368:34375] = '{-71.1927420905, 72.0894386139, 33.8863005777, -54.3444695176, -63.2928637017, 99.7841614149, 8.39293504489, 37.6393093519};
test_label[4296] = '{-71.1927420905};
test_output[4296] = '{170.976903505};
############ END DEBUG ############*/
test_input[34376:34383] = '{32'hc2a19a4f, 32'hc21edea4, 32'hc24ad538, 32'hc1b0d6fa, 32'h427947a4, 32'hc2455022, 32'hc2619b53, 32'hc2342956};
test_label[4297] = '{32'hc1b0d6fa};
test_output[4297] = '{32'h42a8d991};
/*############ DEBUG ############
test_input[34376:34383] = '{-80.8013804708, -39.7174220065, -50.7082214448, -22.1049690731, 62.31996281, -49.3282562883, -56.4016824633, -45.0403683563};
test_label[4297] = '{-22.1049690731};
test_output[4297] = '{84.4249318831};
############ END DEBUG ############*/
test_input[34384:34391] = '{32'hc24e4f34, 32'hc2bf6d2b, 32'hc234868b, 32'hc2a54fdc, 32'h421a1429, 32'hc29be007, 32'h42a8b341, 32'h42b8951a};
test_label[4298] = '{32'hc2a54fdc};
test_output[4298] = '{32'h432ef292};
/*############ DEBUG ############
test_input[34384:34391] = '{-51.5773461032, -95.7132218394, -45.1313879812, -82.6559769061, 38.519688412, -77.9375498702, 84.3501026476, 92.291215217};
test_label[4298] = '{-82.6559769061};
test_output[4298] = '{174.94754787};
############ END DEBUG ############*/
test_input[34392:34399] = '{32'hc2a97d48, 32'hc10b0a9e, 32'h42687859, 32'hc2785d47, 32'h420246f6, 32'hc288d948, 32'hc129475f, 32'hc23c763e};
test_label[4299] = '{32'h42687859};
test_output[4299] = '{32'h2d0d3580};
/*############ DEBUG ############
test_input[34392:34399] = '{-84.7446901885, -8.69009198828, 58.1175269343, -62.0910925608, 32.5692970868, -68.424377233, -10.5799246172, -47.1154717012};
test_label[4299] = '{58.1175269343};
test_output[4299] = '{8.02680144577e-12};
############ END DEBUG ############*/
test_input[34400:34407] = '{32'h41d88c95, 32'hc2256434, 32'hc2142eec, 32'hc215f547, 32'hc297e5dc, 32'hc2332e1b, 32'hc22ee80c, 32'hc26e6c4b};
test_label[4300] = '{32'hc26e6c4b};
test_output[4300] = '{32'h42ad594a};
/*############ DEBUG ############
test_input[34400:34407] = '{27.0686433221, -41.3478542374, -37.0458203404, -37.4895296381, -75.948945511, -44.7950246395, -43.7266095318, -59.6057529558};
test_label[4300] = '{-59.6057529558};
test_output[4300] = '{86.6743962779};
############ END DEBUG ############*/
test_input[34408:34415] = '{32'hc24bcffc, 32'hc1a4980c, 32'h42681557, 32'hc1f7fea4, 32'hc2b45b0d, 32'hc22a65e3, 32'hc1d027a3, 32'h4283d03e};
test_label[4301] = '{32'hc2b45b0d};
test_output[4301] = '{32'h431c15be};
/*############ DEBUG ############
test_input[34408:34415] = '{-50.953109147, -20.5742415471, 58.0208400285, -30.9993357052, -90.1778337966, -42.5994982947, -26.0193544504, 65.9067192132};
test_label[4301] = '{-90.1778337966};
test_output[4301] = '{156.084928955};
############ END DEBUG ############*/
test_input[34416:34423] = '{32'h42a07f57, 32'h4270cb81, 32'hc2c552f6, 32'h418db8ce, 32'h421dbd45, 32'h42839cb9, 32'hc1e27d16, 32'h42b123db};
test_label[4302] = '{32'h421dbd45};
test_output[4302] = '{32'h42448ab1};
/*############ DEBUG ############
test_input[34416:34423] = '{80.2487133872, 60.1987324631, -98.6620336893, 17.7152357278, 39.4348334631, 65.8060952238, -28.311076911, 88.5700327414};
test_label[4302] = '{39.4348334631};
test_output[4302] = '{49.1354425235};
############ END DEBUG ############*/
test_input[34424:34431] = '{32'hc246caf8, 32'h423d0d31, 32'hc27c4d91, 32'hc238d529, 32'h42adabe0, 32'h41eae0d5, 32'h41f8e120, 32'h407dc67b};
test_label[4303] = '{32'hc246caf8};
test_output[4303] = '{32'h430888ae};
/*############ DEBUG ############
test_input[34424:34431] = '{-49.6982124985, 47.2628836744, -63.0757492588, -46.2081658684, 86.8356964244, 29.3597803483, 31.109924659, 3.96523929467};
test_label[4303] = '{-49.6982124985};
test_output[4303] = '{136.533908923};
############ END DEBUG ############*/
test_input[34432:34439] = '{32'h429c9e77, 32'h41d725ad, 32'h42b05315, 32'h40b8c539, 32'h414c9be3, 32'hc13cae16, 32'h418b852a, 32'h42a28a53};
test_label[4304] = '{32'h41d725ad};
test_output[4304] = '{32'h4275146b};
/*############ DEBUG ############
test_input[34432:34439] = '{78.3095042499, 26.8933959456, 88.1622688382, 5.77407520922, 12.7880578793, -11.7925015493, 17.4400210719, 81.2701621384};
test_label[4304] = '{26.8933959456};
test_output[4304] = '{61.2699406955};
############ END DEBUG ############*/
test_input[34440:34447] = '{32'h4103ca6b, 32'hc1f525fe, 32'hc2aba37e, 32'h423bc651, 32'h41670130, 32'hc2c187d6, 32'h42843e26, 32'h424c3d4f};
test_label[4305] = '{32'hc2c187d6};
test_output[4305] = '{32'h4322e2fe};
/*############ DEBUG ############
test_input[34440:34447] = '{8.23691836239, -30.6435509025, -85.8193240302, 46.9436696837, 14.4377901708, -96.7653028817, 66.1213800209, 51.059872565};
test_label[4305] = '{-96.7653028817};
test_output[4305] = '{162.886683195};
############ END DEBUG ############*/
test_input[34448:34455] = '{32'h41d5f9d4, 32'hc28645bd, 32'hc206f150, 32'hc255cdb9, 32'h4267f2e9, 32'hc287071a, 32'h3f83fda3, 32'h409ddf86};
test_label[4306] = '{32'h409ddf86};
test_output[4306] = '{32'h425436f8};
/*############ DEBUG ############
test_input[34448:34455] = '{26.7469872503, -67.1362043407, -33.7356556752, -53.450899554, 57.9872163303, -67.5138691127, 1.03117787837, 4.93353554306};
test_label[4306] = '{4.93353554306};
test_output[4306] = '{53.0536807872};
############ END DEBUG ############*/
test_input[34456:34463] = '{32'hc28cf2d3, 32'h4293d6ce, 32'hc2b24aba, 32'hc2af572b, 32'h41db2647, 32'hc2a49503, 32'h42b21645, 32'hc2b5078c};
test_label[4307] = '{32'hc2b24aba};
test_output[4307] = '{32'h4332307f};
/*############ DEBUG ############
test_input[34456:34463] = '{-70.4742678195, 73.9195405636, -89.1459468007, -87.6702466185, 27.3936894485, -82.2910371732, 89.0434974312, -90.5147381108};
test_label[4307] = '{-89.1459468007};
test_output[4307] = '{178.189444502};
############ END DEBUG ############*/
test_input[34464:34471] = '{32'hc29d4d24, 32'h41145234, 32'h42507b4e, 32'h41f503f9, 32'hbf722f08, 32'h42ad93e8, 32'hc2916b7b, 32'h42b7d126};
test_label[4308] = '{32'h41145234};
test_output[4308] = '{32'h42a549ec};
/*############ DEBUG ############
test_input[34464:34471] = '{-78.6506676925, 9.27006891649, 52.1204131253, 30.6269396521, -0.946030133005, 86.7888777477, -72.7099190783, 91.9084895726};
test_label[4308] = '{9.27006891649};
test_output[4308] = '{82.6443811999};
############ END DEBUG ############*/
test_input[34472:34479] = '{32'h41c2f889, 32'h4271947a, 32'hc2b26518, 32'h4266cb2d, 32'h41933df1, 32'hc2477739, 32'hc2a56eba, 32'hc1a6c066};
test_label[4309] = '{32'h41933df1};
test_output[4309] = '{32'h42283854};
/*############ DEBUG ############
test_input[34472:34479] = '{24.3713559209, 60.3949956194, -89.1974459806, 57.6984147661, 18.4052450475, -49.8664277254, -82.7162605372, -20.8439436707};
test_label[4309] = '{18.4052450475};
test_output[4309] = '{42.0550097941};
############ END DEBUG ############*/
test_input[34480:34487] = '{32'hc15a5aaf, 32'hc29d4cb7, 32'hc232bd75, 32'h42b995c4, 32'hc2bcc096, 32'hc10f6091, 32'h419b75ed, 32'hc00a0cb4};
test_label[4310] = '{32'hc10f6091};
test_output[4310] = '{32'h42cb81d6};
/*############ DEBUG ############
test_input[34480:34487] = '{-13.647139549, -78.6498312067, -44.6850174066, 92.7925119659, -94.3761447401, -8.96107579114, 19.4325809598, -2.15702536331};
test_label[4310] = '{-8.96107579114};
test_output[4310] = '{101.753587757};
############ END DEBUG ############*/
test_input[34488:34495] = '{32'h41b9c9ec, 32'h42c21de0, 32'h416bf729, 32'h42750a54, 32'hc2b527d5, 32'h4288c5b6, 32'h4286c2cd, 32'hc20b128a};
test_label[4311] = '{32'h41b9c9ec};
test_output[4311] = '{32'h4293ab65};
/*############ DEBUG ############
test_input[34488:34495] = '{23.2235941906, 97.0583459308, 14.7478415403, 61.2600856922, -90.5777937018, 68.3861566212, 67.3804722743, -34.768104465};
test_label[4311] = '{23.2235941906};
test_output[4311] = '{73.8347517402};
############ END DEBUG ############*/
test_input[34496:34503] = '{32'hc2c052ae, 32'h423cea2b, 32'hc2148849, 32'hc267e5e4, 32'h41c699a6, 32'h4264e081, 32'h42639082, 32'h423b2c4c};
test_label[4312] = '{32'hc267e5e4};
test_output[4312] = '{32'h42e778f9};
/*############ DEBUG ############
test_input[34496:34503] = '{-96.1614804848, 47.2286802875, -37.1330911312, -57.9745016052, 24.8250231686, 57.2192403115, 56.8911205444, 46.793257461};
test_label[4312] = '{-57.9745016052};
test_output[4312] = '{115.736270972};
############ END DEBUG ############*/
test_input[34504:34511] = '{32'h4124d6cf, 32'h42870df1, 32'h429a66d4, 32'h42784287, 32'h4165d874, 32'hc29b049f, 32'hc2c29c42, 32'h41eb1dff};
test_label[4313] = '{32'h42784287};
test_output[4313] = '{32'h41722cc4};
/*############ DEBUG ############
test_input[34504:34511] = '{10.302443844, 67.5272259545, 77.2008355217, 62.0649693972, 14.365345085, -77.5090268768, -97.3051878359, 29.3896470071};
test_label[4313] = '{62.0649693972};
test_output[4313] = '{15.1359293119};
############ END DEBUG ############*/
test_input[34512:34519] = '{32'hc0a07a2e, 32'hc254e3a5, 32'hc224876a, 32'hc2950b7a, 32'h42c1e82b, 32'h429bd86f, 32'h428af05b, 32'h42c2794d};
test_label[4314] = '{32'h42c1e82b};
test_output[4314] = '{32'h3f584ac3};
/*############ DEBUG ############
test_input[34512:34519] = '{-5.01491438939, -53.2223094668, -41.1322395459, -74.522412751, 96.953452267, 77.9227192468, 69.4694477637, 97.2369181041};
test_label[4314] = '{96.953452267};
test_output[4314] = '{0.844890762557};
############ END DEBUG ############*/
test_input[34520:34527] = '{32'h426bc5e2, 32'hc2630cb0, 32'hc2863cd7, 32'hc2c58147, 32'hc29e82d8, 32'h41ad15b4, 32'h42b3c1e6, 32'h42107bbf};
test_label[4315] = '{32'h41ad15b4};
test_output[4315] = '{32'h42887c79};
/*############ DEBUG ############
test_input[34520:34527] = '{58.9432436064, -56.7623893009, -67.1188253458, -98.752494446, -79.255555843, 21.635596327, 89.8787051068, 36.120844579};
test_label[4315] = '{21.635596327};
test_output[4315] = '{68.2431087798};
############ END DEBUG ############*/
test_input[34528:34535] = '{32'hc123ca88, 32'h429e4c3b, 32'h41ed7800, 32'hc280f79b, 32'hc2b3bc6a, 32'h42131bfc, 32'h41324234, 32'h428fe052};
test_label[4316] = '{32'hc123ca88};
test_output[4316] = '{32'h42b2c5ec};
/*############ DEBUG ############
test_input[34528:34535] = '{-10.236946006, 79.1488838656, 29.6835941277, -64.4836072697, -89.8679994259, 36.7773303155, 11.1411632398, 71.9381277061};
test_label[4316] = '{-10.236946006};
test_output[4316] = '{89.3865681974};
############ END DEBUG ############*/
test_input[34536:34543] = '{32'hc0b867b5, 32'hc1b76110, 32'hc2c5a621, 32'h427d813e, 32'h42b4ed34, 32'hc291fffb, 32'hc2bd4a35, 32'h42ade08c};
test_label[4317] = '{32'h42b4ed34};
test_output[4317] = '{32'h3cedda07};
/*############ DEBUG ############
test_input[34536:34543] = '{-5.76265943798, -22.9223932608, -98.8244694309, 63.376212337, 90.4632850535, -72.9999602934, -94.6449347124, 86.9385713809};
test_label[4317] = '{90.4632850535};
test_output[4317] = '{0.0290346274489};
############ END DEBUG ############*/
test_input[34544:34551] = '{32'hc235b138, 32'hc28e2cca, 32'h419b8317, 32'hc25a4e76, 32'hc18ed8f5, 32'hc298466f, 32'hc245ad11, 32'hc189603c};
test_label[4318] = '{32'hc25a4e76};
test_output[4318] = '{32'h42940801};
/*############ DEBUG ############
test_input[34544:34551] = '{-45.4230647752, -71.0874755621, 19.4390094234, -54.5766235281, -17.8559357246, -76.1375657817, -49.4190118051, -17.1719890597};
test_label[4318] = '{-54.5766235281};
test_output[4318] = '{74.0156329516};
############ END DEBUG ############*/
test_input[34552:34559] = '{32'hc2adfdda, 32'h426929de, 32'hc24d284f, 32'hc2978aa4, 32'h419d5673, 32'h4209afa5, 32'h4131395c, 32'hc134a985};
test_label[4319] = '{32'hc2adfdda};
test_output[4319] = '{32'h43114964};
/*############ DEBUG ############
test_input[34552:34559] = '{-86.9958004666, 58.2908861153, -51.2893635458, -75.7707846185, 19.6672106213, 34.4215290202, 11.0765035513, -11.2913861871};
test_label[4319] = '{-86.9958004666};
test_output[4319] = '{145.286686582};
############ END DEBUG ############*/
test_input[34560:34567] = '{32'h424591a9, 32'hc286a9a4, 32'hc2a2dad5, 32'h420548c7, 32'hc0a8bde1, 32'h4056bc91, 32'hc1bfe8b6, 32'h41dd5f33};
test_label[4320] = '{32'hc1bfe8b6};
test_output[4320] = '{32'h4292c302};
/*############ DEBUG ############
test_input[34560:34567] = '{49.3922456162, -67.3313327346, -81.4274065575, 33.3210724127, -5.27317879295, 3.35525928298, -23.9886292077, 27.6714837857};
test_label[4320] = '{-23.9886292077};
test_output[4320] = '{73.3808749291};
############ END DEBUG ############*/
test_input[34568:34575] = '{32'hc1b0387a, 32'hc20a065b, 32'h4237e616, 32'h4268cce7, 32'hc2aa9eb3, 32'hc21d06ec, 32'hc20d367f, 32'hc0ac6c8a};
test_label[4321] = '{32'hc1b0387a};
test_output[4321] = '{32'h42a07493};
/*############ DEBUG ############
test_input[34568:34575] = '{-22.0275764326, -34.5062049147, 45.9746945609, 58.2001013912, -85.3099557427, -39.2567601064, -35.3032186051, -5.3882493785};
test_label[4321] = '{-22.0275764326};
test_output[4321] = '{80.227682728};
############ END DEBUG ############*/
test_input[34576:34583] = '{32'h4129f381, 32'h4271dd49, 32'h412dba6a, 32'hc1e898f1, 32'hc186151d, 32'h42bf8f55, 32'hc29d1436, 32'h3f30567c};
test_label[4322] = '{32'h4271dd49};
test_output[4322] = '{32'h420d4161};
/*############ DEBUG ############
test_input[34576:34583] = '{10.6219488194, 60.4660996669, 10.8580111214, -29.0746784487, -16.7603092755, 95.7799457871, -78.5394763796, 0.68881962719};
test_label[4322] = '{60.4660996669};
test_output[4322] = '{35.3138461202};
############ END DEBUG ############*/
test_input[34584:34591] = '{32'hc182c698, 32'hc0dbf9d0, 32'hc29a0c52, 32'hc28341bd, 32'hc2c39964, 32'hc2565240, 32'h414702ff, 32'hc20beb5c};
test_label[4323] = '{32'h414702ff};
test_output[4323] = '{32'h318cdba0};
/*############ DEBUG ############
test_input[34584:34591] = '{-16.3469700114, -6.87424470805, -77.0240638082, -65.6283942483, -97.7995901871, -53.5803223564, 12.4382318754, -34.9798420455};
test_label[4323] = '{12.4382318754};
test_output[4323] = '{4.09950463306e-09};
############ END DEBUG ############*/
test_input[34592:34599] = '{32'h42006997, 32'h41d39f12, 32'hc0eaf601, 32'hc24e2022, 32'hc2627175, 32'hc2361be5, 32'hc237f585, 32'h42677f2a};
test_label[4324] = '{32'hc2627175};
test_output[4324] = '{32'h42e4f850};
/*############ DEBUG ############
test_input[34592:34599] = '{32.1031154779, 26.4526702042, -7.34252984967, -51.5313794928, -56.6107997081, -45.5272403542, -45.9897637944, 57.8741834435};
test_label[4324] = '{-56.6107997081};
test_output[4324] = '{114.484983152};
############ END DEBUG ############*/
test_input[34600:34607] = '{32'hc2b0b6d7, 32'hc20b3b0a, 32'hc1749e22, 32'h42140ad8, 32'h42854d3b, 32'h40082e48, 32'h425f847c, 32'h42b5215e};
test_label[4325] = '{32'h425f847c};
test_output[4325] = '{32'h420abe41};
/*############ DEBUG ############
test_input[34600:34607] = '{-88.357110788, -34.807654366, -15.2886063817, 37.010589652, 66.6508396689, 2.12782488922, 55.879378699, 90.565172059};
test_label[4325] = '{55.879378699};
test_output[4325] = '{34.68579336};
############ END DEBUG ############*/
test_input[34608:34615] = '{32'h42413f84, 32'h42691162, 32'h4294429d, 32'h41438f3a, 32'h42945f06, 32'h4202f9eb, 32'h42787649, 32'h42468ff2};
test_label[4326] = '{32'h42413f84};
test_output[4326] = '{32'h41d4509a};
/*############ DEBUG ############
test_input[34608:34615] = '{48.3120263142, 58.2669770265, 74.1301044843, 12.2224678224, 74.1855903859, 32.7440590215, 62.1155143316, 49.6405700028};
test_label[4326] = '{48.3120263142};
test_output[4326] = '{26.5393560941};
############ END DEBUG ############*/
test_input[34616:34623] = '{32'hc286fc4b, 32'hc2338ac5, 32'h41b44af8, 32'hc29de300, 32'hbf0ac407, 32'h42259351, 32'h4212832d, 32'hc2bf4b39};
test_label[4327] = '{32'hbf0ac407};
test_output[4327] = '{32'h4227c710};
/*############ DEBUG ############
test_input[34616:34623] = '{-67.4927569908, -44.8855155428, 22.5366067859, -78.9433591209, -0.542053627294, 41.393863281, 36.6281021651, -95.6469218905};
test_label[4327] = '{-0.542053627294};
test_output[4327] = '{41.9443972585};
############ END DEBUG ############*/
test_input[34624:34631] = '{32'hc2163be1, 32'h42a23dc1, 32'h429e547d, 32'h4290f8cc, 32'hc2ab42f5, 32'h42c5bf74, 32'h41b8a30b, 32'h42c3121d};
test_label[4328] = '{32'h42c3121d};
test_output[4328] = '{32'h3fc924b4};
/*############ DEBUG ############
test_input[34624:34631] = '{-37.5584760003, 81.1206126672, 79.1650189863, 72.4859311113, -85.6307743856, 98.873935441, 23.0796102288, 97.5353777558};
test_label[4328] = '{97.5353777558};
test_output[4328] = '{1.57143263425};
############ END DEBUG ############*/
test_input[34632:34639] = '{32'hc2943606, 32'h41475fd7, 32'h4215c397, 32'h41b2bfd5, 32'hc1b44585, 32'h4257d022, 32'hbeec8343, 32'h42847e08};
test_label[4329] = '{32'h4257d022};
test_output[4329] = '{32'h4144afbc};
/*############ DEBUG ############
test_input[34632:34639] = '{-74.1055170895, 12.4608986987, 37.441006845, 22.3436688, -22.5339454945, 53.9532542231, -0.461938947563, 66.2461534736};
test_label[4329] = '{53.9532542231};
test_output[4329] = '{12.2929038347};
############ END DEBUG ############*/
test_input[34640:34647] = '{32'hc20ea323, 32'hc1909afd, 32'h4252ce9f, 32'h42b0ed66, 32'hc26e4030, 32'hc13203c9, 32'h4248c645, 32'h4281e5af};
test_label[4330] = '{32'h42b0ed66};
test_output[4330] = '{32'h2e86d310};
/*############ DEBUG ############
test_input[34640:34647] = '{-35.6593114326, -18.0756782761, 52.7017787319, 88.4636651459, -59.5626816844, -11.1259239682, 50.193621828, 64.9486000585};
test_label[4330] = '{88.4636651459};
test_output[4330] = '{6.13110673361e-11};
############ END DEBUG ############*/
test_input[34648:34655] = '{32'h4106c9cd, 32'h41960476, 32'hc102e556, 32'hbf9a42b8, 32'hc22902f3, 32'h42a19298, 32'hc28935fe, 32'h3f4f1e42};
test_label[4331] = '{32'hbf9a42b8};
test_output[4331] = '{32'h42a3fba2};
/*############ DEBUG ############
test_input[34648:34655] = '{8.42426793833, 18.7521776438, -8.1809897455, -1.20516111962, -42.2528807083, 80.7863121508, -68.6054510068, 0.809055429293};
test_label[4331] = '{-1.20516111962};
test_output[4331] = '{81.9914732705};
############ END DEBUG ############*/
test_input[34656:34663] = '{32'h400b7db3, 32'h414b91d0, 32'h4222b6c1, 32'hc2945c99, 32'hc001617d, 32'h402afe12, 32'hc1b8b81a, 32'h4291f16b};
test_label[4332] = '{32'h402afe12};
test_output[4332] = '{32'h428c997b};
/*############ DEBUG ############
test_input[34656:34663] = '{2.1795470959, 12.72309866, 40.6784718605, -74.180853756, -2.02157523282, 2.67175716424, -23.089893506, 72.9715228512};
test_label[4332] = '{2.67175716424};
test_output[4332] = '{70.2997656869};
############ END DEBUG ############*/
test_input[34664:34671] = '{32'hc21f402c, 32'h4275f1fe, 32'h41d75b34, 32'h41af07c1, 32'hc22733aa, 32'hc1dd328d, 32'hc25f20d0, 32'hc21fed7e};
test_label[4333] = '{32'hc21f402c};
test_output[4333] = '{32'h42ca9915};
/*############ DEBUG ############
test_input[34664:34671] = '{-39.8126679144, 61.4863196824, 26.919532761, 21.8787869024, -41.8004530093, -27.6496821108, -55.7820441393, -39.9819256412};
test_label[4333] = '{-39.8126679144};
test_output[4333] = '{101.298987597};
############ END DEBUG ############*/
test_input[34672:34679] = '{32'hc299eb60, 32'hc1c6334b, 32'hc1ec9695, 32'h424c649b, 32'hc29448a0, 32'h428b7118, 32'hc167e785, 32'h42c7aba7};
test_label[4334] = '{32'hc1ec9695};
test_output[4334] = '{32'h430168a6};
/*############ DEBUG ############
test_input[34672:34679] = '{-76.959716008, -24.7750455261, -29.5735270972, 51.0982461923, -74.1418470678, 69.7208836302, -14.494023564, 99.8352584411};
test_label[4334] = '{-29.5735270972};
test_output[4334] = '{129.408785538};
############ END DEBUG ############*/
test_input[34680:34687] = '{32'hc280aa23, 32'h4246eb44, 32'hc273379c, 32'hc2beb75b, 32'h429c188f, 32'hc17d2323, 32'hc28dcbae, 32'hc176bb69};
test_label[4335] = '{32'hc176bb69};
test_output[4335] = '{32'h42baeffc};
/*############ DEBUG ############
test_input[34680:34687] = '{-64.3323017585, 49.729752381, -60.8043065301, -95.3581195152, 78.0479673293, -15.8210782908, -70.8978131695, -15.4207541465};
test_label[4335] = '{-15.4207541465};
test_output[4335] = '{93.4687214758};
############ END DEBUG ############*/
test_input[34688:34695] = '{32'hbfed6089, 32'h41388960, 32'h42827f63, 32'h42a7e657, 32'hc25be37d, 32'hc24517db, 32'hc2b21c71, 32'h422b4585};
test_label[4336] = '{32'hc2b21c71};
test_output[4336] = '{32'h432d0164};
/*############ DEBUG ############
test_input[34688:34695] = '{-1.85450848622, 11.5335386464, 65.2488058802, 83.9498827471, -54.9721578813, -49.273295597, -89.0555520128, 42.817888292};
test_label[4336] = '{-89.0555520128};
test_output[4336] = '{173.005434767};
############ END DEBUG ############*/
test_input[34696:34703] = '{32'h41806e39, 32'hc29a2631, 32'h420a0825, 32'hc2bf2c1d, 32'hc28d3061, 32'h429d4a5a, 32'hc2c52ee7, 32'h42656117};
test_label[4337] = '{32'hc29a2631};
test_output[4337] = '{32'h431bb845};
/*############ DEBUG ############
test_input[34696:34703] = '{16.0538199341, -77.0745901042, 34.5079549114, -95.5861574754, -70.5944879512, 78.6452181954, -98.5916081707, 57.3448139564};
test_label[4337] = '{-77.0745901042};
test_output[4337] = '{155.7198083};
############ END DEBUG ############*/
test_input[34704:34711] = '{32'hc28d12af, 32'h40e6a672, 32'hc2652d97, 32'h425cf460, 32'h429a17e1, 32'h40ed6143, 32'hc1277c8a, 32'hc1ebc88e};
test_label[4338] = '{32'h425cf460};
test_output[4338] = '{32'h41ae76c2};
/*############ DEBUG ############
test_input[34704:34711] = '{-70.5364916867, 7.20781815669, -57.2945227068, 55.2386485868, 77.0466362468, 7.41812287966, -10.4679049416, -29.4729264565};
test_label[4338] = '{55.2386485868};
test_output[4338] = '{21.8079876604};
############ END DEBUG ############*/
test_input[34712:34719] = '{32'h3e81acfa, 32'h4291e98c, 32'h41ed2066, 32'h4229fdaf, 32'h411c36fc, 32'hc2b56d05, 32'h42b0ad1f, 32'hc24dd6e5};
test_label[4339] = '{32'h42b0ad1f};
test_output[4339] = '{32'h34602cef};
/*############ DEBUG ############
test_input[34712:34719] = '{0.253272834121, 72.9561448097, 29.6408201182, 42.4977367544, 9.76342413112, -90.712927048, 88.338130815, -51.4598584814};
test_label[4339] = '{88.338130815};
test_output[4339] = '{2.08779720546e-07};
############ END DEBUG ############*/
test_input[34720:34727] = '{32'h41b99f4d, 32'h4296e350, 32'hc2ba0e16, 32'hc2a9b37b, 32'hc2bc7eb5, 32'hc26346e1, 32'h41d77aea, 32'h423f87e7};
test_label[4340] = '{32'h4296e350};
test_output[4340] = '{32'h2b96e800};
/*############ DEBUG ############
test_input[34720:34727] = '{23.2027827587, 75.4439724902, -93.0275139936, -84.8505508359, -94.2474782672, -56.8192193283, 26.9350157055, 47.8827181303};
test_label[4340] = '{75.4439724902};
test_output[4340] = '{1.07225339718e-12};
############ END DEBUG ############*/
test_input[34728:34735] = '{32'hc29004e5, 32'hc0d08323, 32'hc2a7fc9d, 32'h3d057c0b, 32'h421aa210, 32'hc114f15e, 32'hc18c4445, 32'hc1c95a27};
test_label[4341] = '{32'hc1c95a27};
test_output[4341] = '{32'h427f4f23};
/*############ DEBUG ############
test_input[34728:34735] = '{-72.0095573464, -6.51600774745, -83.9933856537, 0.0325889984655, 38.6582636657, -9.30892725839, -17.533335031, -25.1690187691};
test_label[4341] = '{-25.1690187691};
test_output[4341] = '{63.8272824348};
############ END DEBUG ############*/
test_input[34736:34743] = '{32'h429959ed, 32'hc2ac4876, 32'h4239df35, 32'hc25cda5f, 32'hc237d8c2, 32'h4284f6f5, 32'h40202a23, 32'hc2919459};
test_label[4342] = '{32'hc2919459};
test_output[4342] = '{32'h43157725};
/*############ DEBUG ############
test_input[34736:34743] = '{76.6756336745, -86.1415288659, 46.4679771821, -55.2132535721, -45.96167941, 66.4823400933, 2.50257175079, -72.7897428612};
test_label[4342] = '{-72.7897428612};
test_output[4342] = '{149.465413955};
############ END DEBUG ############*/
test_input[34744:34751] = '{32'h4233ff6b, 32'h41dc2944, 32'h4284cbd2, 32'hc11ac073, 32'h41d5367d, 32'hc29f19db, 32'hc25d0568, 32'hc2bca251};
test_label[4343] = '{32'hc2bca251};
test_output[4343] = '{32'h4320b712};
/*############ DEBUG ############
test_input[34744:34751] = '{44.9994316727, 27.5201482963, 66.3980888845, -9.67198483025, 26.6516052981, -79.5504954402, -55.2552785872, -94.3170271754};
test_label[4343] = '{-94.3170271754};
test_output[4343] = '{160.71511606};
############ END DEBUG ############*/
test_input[34752:34759] = '{32'h4296189c, 32'h428d5dd8, 32'h4169c2eb, 32'h422ba228, 32'h41c3de10, 32'hc237eae8, 32'h42b84488, 32'hc207b7e8};
test_label[4344] = '{32'h4296189c};
test_output[4344] = '{32'h4188afb1};
/*############ DEBUG ############
test_input[34752:34759] = '{75.0480614289, 70.6832918389, 14.6100871139, 42.9083568972, 24.4834284471, -45.9794010936, 92.1338489742, -33.9295956432};
test_label[4344] = '{75.0480614289};
test_output[4344] = '{17.0857875838};
############ END DEBUG ############*/
test_input[34760:34767] = '{32'hc1857fc3, 32'h415686fc, 32'h428c56da, 32'hc2b0a4da, 32'h42a48b17, 32'h41caa796, 32'h421c7c24, 32'h42461e9a};
test_label[4345] = '{32'h42461e9a};
test_output[4345] = '{32'h4202f795};
/*############ DEBUG ############
test_input[34760:34767] = '{-16.6873834617, 13.4079549264, 70.1696322834, -88.3219737378, 82.2716577104, 25.3318286453, 39.1212314894, 49.5298832255};
test_label[4345] = '{49.5298832255};
test_output[4345] = '{32.7417800331};
############ END DEBUG ############*/
test_input[34768:34775] = '{32'hc2a82a5b, 32'h406afa2b, 32'h4165c55c, 32'hc153833c, 32'h42c542a1, 32'hc15ea5af, 32'hc2a1d884, 32'hc1bed9e8};
test_label[4346] = '{32'hc15ea5af};
test_output[4346] = '{32'h42e11757};
/*############ DEBUG ############
test_input[34768:34775] = '{-84.0827248947, 3.67151899796, 14.3606835272, -13.2195399775, 98.6301321093, -13.9154501532, -80.9228847162, -23.85639915};
test_label[4346] = '{-13.9154501532};
test_output[4346] = '{112.545582263};
############ END DEBUG ############*/
test_input[34776:34783] = '{32'hc213a516, 32'h4154458f, 32'hc2c6f0dc, 32'h428bc49f, 32'hc26fdeb4, 32'hc2b0cd69, 32'h42c6f9db, 32'h42b1340a};
test_label[4347] = '{32'hc2c6f0dc};
test_output[4347] = '{32'h4346f55c};
/*############ DEBUG ############
test_input[34776:34783] = '{-36.9112151326, 13.2669824533, -99.4704247436, 69.8840271189, -59.9674830147, -88.4011941896, 99.487998892, 88.6016417739};
test_label[4347] = '{-99.4704247436};
test_output[4347] = '{198.958442347};
############ END DEBUG ############*/
test_input[34784:34791] = '{32'hc2b2ee41, 32'h40e1c4e0, 32'h427b0ce3, 32'hc04de2ff, 32'h42111b4c, 32'hc2a99cdb, 32'h3ec634f2, 32'hc232ad1f};
test_label[4348] = '{32'h40e1c4e0};
test_output[4348] = '{32'h425ed447};
/*############ DEBUG ############
test_input[34784:34791] = '{-89.465338646, 7.05528266817, 62.7625853042, -3.21697976787, 36.2766552605, -84.8063562959, 0.387122703775, -44.6690625006};
test_label[4348] = '{7.05528266817};
test_output[4348] = '{55.7073026361};
############ END DEBUG ############*/
test_input[34792:34799] = '{32'hc1d06356, 32'h41f4da2e, 32'h42baaff0, 32'h41c71809, 32'h423207c6, 32'h42157a28, 32'h427be1b8, 32'h41c3e246};
test_label[4349] = '{32'h42157a28};
test_output[4349] = '{32'h425fe5b8};
/*############ DEBUG ############
test_input[34792:34799] = '{-26.0485038571, 30.6065332624, 93.3436284495, 24.8867367968, 44.5075911928, 37.3692928642, 62.9704300317, 24.4854855381};
test_label[4349] = '{37.3692928642};
test_output[4349] = '{55.9743355853};
############ END DEBUG ############*/
test_input[34800:34807] = '{32'h42a72d79, 32'h42b993fd, 32'hc124eb39, 32'h40b11dd4, 32'hc259b4f4, 32'h427196f6, 32'h4145bb2d, 32'hc2a3818a};
test_label[4350] = '{32'hc259b4f4};
test_output[4350] = '{32'h43133742};
/*############ DEBUG ############
test_input[34800:34807] = '{83.588810713, 92.789038177, -10.3074270228, 5.53489098836, -54.4267134974, 60.3974233623, 12.3581970415, -81.7530049402};
test_label[4350] = '{-54.4267134974};
test_output[4350] = '{147.215852686};
############ END DEBUG ############*/
test_input[34808:34815] = '{32'hc281fe1e, 32'hc251bc71, 32'hc2264022, 32'h4280fa7b, 32'h4227fcfe, 32'h4256d2c0, 32'h42a4309c, 32'h4176ae04};
test_label[4351] = '{32'h42a4309c};
test_output[4351] = '{32'h32c20f05};
/*############ DEBUG ############
test_input[34808:34815] = '{-64.9963225103, -52.4340236746, -41.5626284109, 64.4892203343, 41.9970636503, 53.7058103662, 82.0949374992, 15.4174841409};
test_label[4351] = '{82.0949374992};
test_output[4351] = '{2.25914022265e-08};
############ END DEBUG ############*/
test_input[34816:34823] = '{32'hc1892e39, 32'hc22b692e, 32'hc28254aa, 32'h4220db6d, 32'h411380e9, 32'hc1864ee7, 32'h41e29a22, 32'h429f9dad};
test_label[4352] = '{32'h4220db6d};
test_output[4352] = '{32'h421e5fed};
/*############ DEBUG ############
test_input[34816:34823] = '{-17.1475687814, -42.85271294, -65.1653579937, 40.2142841426, 9.21897177829, -16.7885274055, 28.3252609379, 79.8079629974};
test_label[4352] = '{40.2142841426};
test_output[4352] = '{39.5936788548};
############ END DEBUG ############*/
test_input[34824:34831] = '{32'h42934156, 32'hc1cad99f, 32'h41970740, 32'hc2068913, 32'h429f6c53, 32'hc1bbfef6, 32'h420f8704, 32'hc1ede2d2};
test_label[4353] = '{32'hc1cad99f};
test_output[4353] = '{32'h42d223e5};
/*############ DEBUG ############
test_input[34824:34831] = '{73.6276130051, -25.3562595623, 18.8785397908, -33.6338624303, 79.7115682218, -23.4994924744, 35.8818501436, -29.7357519515};
test_label[4353] = '{-25.3562595623};
test_output[4353] = '{105.070104335};
############ END DEBUG ############*/
test_input[34832:34839] = '{32'hc133d6bc, 32'h424b842b, 32'hc2b15da6, 32'hc1b8b966, 32'hc1be9ec6, 32'hc2c03f72, 32'h4223e490, 32'h41c8fc11};
test_label[4354] = '{32'hc133d6bc};
test_output[4354] = '{32'h427879e7};
/*############ DEBUG ############
test_input[34832:34839] = '{-11.2399253492, 50.8790704829, -88.6829074235, -23.0905264421, -23.8275260863, -96.123917618, 40.9732070955, 25.1230789264};
test_label[4354] = '{-11.2399253492};
test_output[4354] = '{62.1190457122};
############ END DEBUG ############*/
test_input[34840:34847] = '{32'hc2aeece1, 32'hc1f6d6f5, 32'hc1e4d2de, 32'hc24003e0, 32'hc2a7912d, 32'h424e9e7b, 32'hc24e6fa0, 32'hbf93b278};
test_label[4355] = '{32'hc24003e0};
test_output[4355] = '{32'h42c7512d};
/*############ DEBUG ############
test_input[34840:34847] = '{-87.4626575871, -30.8549594035, -28.6029622093, -48.0037824021, -83.7835446708, 51.6547675493, -51.6090097754, -1.15388393047};
test_label[4355] = '{-48.0037824021};
test_output[4355] = '{99.6585499513};
############ END DEBUG ############*/
test_input[34848:34855] = '{32'hc1d66009, 32'h428191c8, 32'h41966f95, 32'h40f57d2d, 32'h42803fe6, 32'h4173f9e1, 32'h403717f8, 32'h40e37307};
test_label[4356] = '{32'h41966f95};
test_output[4356] = '{32'h4239966f};
/*############ DEBUG ############
test_input[34848:34855] = '{-26.7968913572, 64.7847296504, 18.8044833825, 7.671530431, 64.1247990988, 15.2485052977, 2.86083787441, 7.10779163827};
test_label[4356] = '{18.8044833825};
test_output[4356] = '{46.3969066282};
############ END DEBUG ############*/
test_input[34856:34863] = '{32'hc13361fa, 32'hc28227c7, 32'h42a295cf, 32'h4285c7f5, 32'hc2a21efd, 32'hc29de38a, 32'h42311c2b, 32'hc17bb0eb};
test_label[4357] = '{32'h4285c7f5};
test_output[4357] = '{32'h41666ed0};
/*############ DEBUG ############
test_input[34856:34863] = '{-11.211420323, -65.0776934372, 81.2925945709, 66.8905414933, -81.0605246596, -78.9444101714, 44.2775077408, -15.7306930213};
test_label[4357] = '{66.8905414933};
test_output[4357] = '{14.4020536338};
############ END DEBUG ############*/
test_input[34864:34871] = '{32'hc1a7283a, 32'h41b6ee0b, 32'h41023e84, 32'h424a88f6, 32'hc2913767, 32'h42212b5c, 32'h418a20d6, 32'hc0443fd8};
test_label[4358] = '{32'hc1a7283a};
test_output[4358] = '{32'h428f0e8d};
/*############ DEBUG ############
test_input[34864:34871] = '{-20.8946415992, 22.8662315186, 8.14026214038, 50.6337490742, -72.6082085571, 40.2923416983, 17.266034089, -3.06639665903};
test_label[4358] = '{-20.8946415992};
test_output[4358] = '{71.5284229417};
############ END DEBUG ############*/
test_input[34872:34879] = '{32'hc10874f4, 32'h41e2f681, 32'hc18c4442, 32'hc0a27198, 32'hc1994acd, 32'hc0af98da, 32'h42665fab, 32'hc29ca05c};
test_label[4359] = '{32'hc1994acd};
test_output[4359] = '{32'h42998289};
/*############ DEBUG ############
test_input[34872:34879] = '{-8.52855346316, 28.370363211, -17.5333286499, -5.07636646352, -19.1615247017, -5.48740848038, 57.5934251231, -78.3132039304};
test_label[4359] = '{-19.1615247017};
test_output[4359] = '{76.7549498248};
############ END DEBUG ############*/
test_input[34880:34887] = '{32'h42a51283, 32'hc28b9280, 32'hc215b18c, 32'h42b1e1f7, 32'hc266023a, 32'h4103e7bb, 32'h42a58900, 32'hc2462464};
test_label[4360] = '{32'hc215b18c};
test_output[4360] = '{32'h42fcbca5};
/*############ DEBUG ############
test_input[34880:34887] = '{82.5361572927, -69.7861323897, -37.4233840755, 88.9413356532, -57.5021744583, 8.24407493069, 82.7675801965, -49.5355371978};
test_label[4360] = '{-37.4233840755};
test_output[4360] = '{126.368449138};
############ END DEBUG ############*/
test_input[34888:34895] = '{32'h41d29259, 32'hc2146277, 32'hc1025fda, 32'hc28a333d, 32'h42790336, 32'hbfcabee9, 32'h410db64b, 32'h427fc678};
test_label[4361] = '{32'h427fc678};
test_output[4361] = '{32'h3e2d4af7};
/*############ DEBUG ############
test_input[34888:34895] = '{26.3214592887, -37.0961578696, -8.14840129415, -69.1000717983, 62.2531358641, -1.58395114676, 8.85700550969, 63.9438161849};
test_label[4361] = '{63.9438161849};
test_output[4361] = '{0.169231280264};
############ END DEBUG ############*/
test_input[34896:34903] = '{32'hc1f1d9b4, 32'hbfc48594, 32'hc2101d38, 32'h42b72092, 32'hc2a817d9, 32'h42b101f5, 32'h40efced0, 32'h4094ab5c};
test_label[4362] = '{32'h42b101f5};
test_output[4362] = '{32'h4046c279};
/*############ DEBUG ############
test_input[34896:34903] = '{-30.2312994894, -1.53532642221, -36.0285328255, 91.5636126105, -84.0465749542, 88.503824109, 7.49399544784, 4.64591800119};
test_label[4362] = '{88.503824109};
test_output[4362] = '{3.10561963766};
############ END DEBUG ############*/
test_input[34904:34911] = '{32'h40aa68d2, 32'hc24f00eb, 32'hc1746119, 32'hc2944342, 32'hc263fece, 32'hc29ce6d8, 32'h40c17c17, 32'h42baa4a1};
test_label[4363] = '{32'hc1746119};
test_output[4363] = '{32'h42d930c4};
/*############ DEBUG ############
test_input[34904:34911] = '{5.32529547651, -51.750896786, -15.2737056026, -74.1313646744, -56.9988336942, -78.4508704584, 6.04639758553, 93.3215386235};
test_label[4363] = '{-15.2737056026};
test_output[4363] = '{108.595244226};
############ END DEBUG ############*/
test_input[34912:34919] = '{32'h41042df8, 32'hc26840e7, 32'hc026eda1, 32'h4245a233, 32'hc1ad137f, 32'hc1c0bc97, 32'hc2266cef, 32'h425c813a};
test_label[4364] = '{32'h4245a233};
test_output[4364] = '{32'h40b71314};
/*############ DEBUG ############
test_input[34912:34919] = '{8.26122249786, -58.0633821581, -2.60825369302, 49.4083984043, -21.6345189354, -24.0920853623, -41.6063811949, 55.1261959334};
test_label[4364] = '{49.4083984043};
test_output[4364] = '{5.7210790813};
############ END DEBUG ############*/
test_input[34920:34927] = '{32'h40dfa274, 32'hc00cbdbc, 32'h4195cde7, 32'h42218beb, 32'h4255e1ef, 32'h426a91b9, 32'hc29c6004, 32'hc26ff45e};
test_label[4365] = '{32'h4255e1ef};
test_output[4365] = '{32'h40a5acad};
/*############ DEBUG ############
test_input[34920:34927] = '{6.98858083799, -2.1990804404, 18.7255385188, 40.3866370968, 53.4706377947, 58.6423072156, -78.187531857, -59.9886414699};
test_label[4365] = '{53.4706377947};
test_output[4365] = '{5.17732847684};
############ END DEBUG ############*/
test_input[34928:34935] = '{32'h42c1e4dd, 32'hc2702d47, 32'hc1dbf44b, 32'hc2bcd1bf, 32'hc2747495, 32'hc25b719b, 32'h4195e5c3, 32'h42a3bdbf};
test_label[4366] = '{32'hc2bcd1bf};
test_output[4366] = '{32'h433f5b4e};
/*############ DEBUG ############
test_input[34928:34935] = '{96.9469965109, -60.0442152196, -27.4942842732, -94.4096618378, -61.1138487725, -54.8609440132, 18.7371883187, 81.8705950889};
test_label[4366] = '{-94.4096618378};
test_output[4366] = '{191.356658632};
############ END DEBUG ############*/
test_input[34936:34943] = '{32'h428eac8b, 32'h417e6db3, 32'hc1a3b783, 32'h42c5d63e, 32'h42c7520e, 32'hc1ee61e5, 32'h42b9c8b4, 32'hc29dbac4};
test_label[4367] = '{32'h42c7520e};
test_output[4367] = '{32'h3ec7d304};
/*############ DEBUG ############
test_input[34936:34943] = '{71.3370005058, 15.9017816216, -20.4646047681, 98.9184438155, 99.6602616441, -29.7978001795, 92.8919958115, -78.8647738186};
test_label[4367] = '{99.6602616441};
test_output[4367] = '{0.390281808795};
############ END DEBUG ############*/
test_input[34944:34951] = '{32'hbf906840, 32'hc232e34a, 32'h4285a54e, 32'hc29bf971, 32'hc20eb0d2, 32'hc21a92b0, 32'h424b5c13, 32'hc287989d};
test_label[4368] = '{32'hc29bf971};
test_output[4368] = '{32'h4310cf60};
/*############ DEBUG ############
test_input[34944:34951] = '{-1.12818149875, -44.7219618978, 66.8228597931, -77.9871935703, -35.6726754412, -38.6432490585, 50.8399162761, -67.7980751451};
test_label[4368] = '{-77.9871935703};
test_output[4368] = '{144.810053478};
############ END DEBUG ############*/
test_input[34952:34959] = '{32'hc2a9fbfe, 32'h418a1f0a, 32'h41ad2a37, 32'h429b3084, 32'hc0883657, 32'h41fc8e1d, 32'h428a1481, 32'hc275e8dc};
test_label[4369] = '{32'h41ad2a37};
test_output[4369] = '{32'h425fcc20};
/*############ DEBUG ############
test_input[34952:34959] = '{-84.9921697519, 17.2651556758, 21.6456126475, 77.5947608777, -4.25663343148, 31.5693914719, 69.0400504635, -61.4774023074};
test_label[4369] = '{21.6456126475};
test_output[4369] = '{55.9493408473};
############ END DEBUG ############*/
test_input[34960:34967] = '{32'h42b373a2, 32'hc03c7602, 32'h41003736, 32'hc29a486b, 32'h42075b68, 32'h427168f3, 32'h42798b0a, 32'h42c27a5f};
test_label[4370] = '{32'h42c27a5f};
test_output[4370] = '{32'h3a0f0d74};
/*############ DEBUG ############
test_input[34960:34967] = '{89.7258427754, -2.94470269454, 8.01347881746, -77.1414430135, 33.8392639141, 60.3524878827, 62.3857811479, 97.2390070996};
test_label[4370] = '{97.2390070996};
test_output[4370] = '{0.000545702180654};
############ END DEBUG ############*/
test_input[34968:34975] = '{32'h42ba76a2, 32'h423e334c, 32'h412f5456, 32'h4264e952, 32'h422439f6, 32'h4254daa9, 32'hc1bb987b, 32'h429a304e};
test_label[4371] = '{32'h412f5456};
test_output[4371] = '{32'h42a48c17};
/*############ DEBUG ############
test_input[34968:34975] = '{93.2317039782, 47.5500944886, 10.9580897282, 57.2278507692, 41.0566029361, 53.2135354565, -23.4494525649, 77.0943451181};
test_label[4371] = '{10.9580897282};
test_output[4371] = '{82.2736143481};
############ END DEBUG ############*/
test_input[34976:34983] = '{32'hc2ad5e04, 32'hc2646b9c, 32'h42a89d10, 32'hc1beb2f8, 32'h41fc56e7, 32'h42c3beb6, 32'hc167d377, 32'h409eb9f1};
test_label[4372] = '{32'hc1beb2f8};
test_output[4372] = '{32'h42f36b74};
/*############ DEBUG ############
test_input[34976:34983] = '{-86.6836208171, -57.1050879235, 84.3067600025, -23.8373866178, 31.5424321333, 97.872484808, -14.4891272351, 4.96019784872};
test_label[4372] = '{-23.8373866178};
test_output[4372] = '{121.709872709};
############ END DEBUG ############*/
test_input[34984:34991] = '{32'hc27e38f6, 32'h4287f92f, 32'h40e3e1ba, 32'h415a69da, 32'h4271f571, 32'hc22c9ddb, 32'hc273b4b5, 32'h41e9c719};
test_label[4373] = '{32'hc27e38f6};
test_output[4373] = '{32'h43038af9};
/*############ DEBUG ############
test_input[34984:34991] = '{-63.5556249925, 67.9866845172, 7.12130430422, 13.6508422681, 60.48968728, -43.1541561253, -60.9264733378, 29.2222148316};
test_label[4373] = '{-63.5556249925};
test_output[4373] = '{131.542864104};
############ END DEBUG ############*/
test_input[34992:34999] = '{32'hc266d8d5, 32'h4216ad03, 32'h41fd647c, 32'hc0f56dad, 32'h428f49e5, 32'hc2584404, 32'h424909ce, 32'h4237f8ee};
test_label[4374] = '{32'hc0f56dad};
test_output[4374] = '{32'h429ea0c0};
/*############ DEBUG ############
test_input[34992:34999] = '{-57.7117516881, 37.6689573202, 31.6740639548, -7.66963792238, 71.6443284407, -54.0664228995, 50.2595751537, 45.9930972167};
test_label[4374] = '{-7.66963792238};
test_output[4374] = '{79.3139663636};
############ END DEBUG ############*/
test_input[35000:35007] = '{32'h42affe87, 32'h419d8f8f, 32'hc015179e, 32'hc1cf78bf, 32'h413494d4, 32'hc2c1bb91, 32'h42a7b703, 32'h405d3ac7};
test_label[4375] = '{32'h413494d4};
test_output[4375] = '{32'h42997404};
/*############ DEBUG ############
test_input[35000:35007] = '{87.9971221588, 19.6950977393, -2.32956644427, -25.9339588647, 11.2863350494, -96.8663369875, 83.8574483039, 3.45671252247};
test_label[4375] = '{11.2863350494};
test_output[4375] = '{76.7265896347};
############ END DEBUG ############*/
test_input[35008:35015] = '{32'h41ce4933, 32'h4263e2cc, 32'h412b66f1, 32'hc24b132e, 32'h41ef3cc1, 32'hc1fee771, 32'h42c11621, 32'hc2833dfc};
test_label[4376] = '{32'h41ef3cc1};
test_output[4376] = '{32'h428546f1};
/*############ DEBUG ############
test_input[35008:35015] = '{25.7857411912, 56.971481785, 10.7126321315, -50.7687309441, 29.9046642297, -31.8630088805, 96.5432210896, -65.6210646464};
test_label[4376] = '{29.9046642297};
test_output[4376] = '{66.6385568599};
############ END DEBUG ############*/
test_input[35016:35023] = '{32'hc0a908cb, 32'hc254851e, 32'hc2ae2ee1, 32'hc21e239f, 32'h41bc7a56, 32'h4172068f, 32'h426b3de6, 32'hc1d50f8a};
test_label[4377] = '{32'h426b3de6};
test_output[4377] = '{32'h26000000};
/*############ DEBUG ############
test_input[35016:35023] = '{-5.28232325224, -53.1299973273, -87.0915622633, -39.5347856224, 23.5597338466, 15.1266015618, 58.8104471707, -26.632587778};
test_label[4377] = '{58.8104471707};
test_output[4377] = '{4.4408920985e-16};
############ END DEBUG ############*/
test_input[35024:35031] = '{32'h4142ba17, 32'h42674f1c, 32'hc28ff167, 32'h427fc633, 32'hc262c5a5, 32'h4245161b, 32'h42065fcc, 32'hc288868e};
test_label[4378] = '{32'h4245161b};
test_output[4378] = '{32'h416ac967};
/*############ DEBUG ############
test_input[35024:35031] = '{12.1704325351, 57.8272553171, -71.9714872021, 63.9435527538, -56.6930124212, 49.2715866007, 33.5935517635, -68.2627998741};
test_label[4378] = '{49.2715866007};
test_output[4378] = '{14.6741707568};
############ END DEBUG ############*/
test_input[35032:35039] = '{32'h4178e963, 32'h42aa882b, 32'hc29d8326, 32'hc2b06e90, 32'h4218b613, 32'h421af1ac, 32'hc22e569b, 32'hc26c41b0};
test_label[4379] = '{32'hc2b06e90};
test_output[4379] = '{32'h432d7b5e};
/*############ DEBUG ############
test_input[35032:35039] = '{15.5569789835, 85.2659553965, -78.7561501122, -88.2159460546, 38.1778051568, 38.7360093443, -43.5845748625, -59.0641460939};
test_label[4379] = '{-88.2159460546};
test_output[4379] = '{173.481901451};
############ END DEBUG ############*/
test_input[35040:35047] = '{32'hc2c371c0, 32'h42852a4a, 32'h42b7b264, 32'hc202272f, 32'h4253ce63, 32'hc26eaa0f, 32'hc293d098, 32'h424f34b6};
test_label[4380] = '{32'hc293d098};
test_output[4380] = '{32'h4325c17e};
/*############ DEBUG ############
test_input[35040:35047] = '{-97.7221699881, 66.5825953373, 91.8484215768, -32.5382635008, 52.9515510537, -59.6660726509, -73.9074073429, 51.8014753482};
test_label[4380] = '{-73.9074073429};
test_output[4380] = '{165.75582892};
############ END DEBUG ############*/
test_input[35048:35055] = '{32'h42187f00, 32'h41e94ed3, 32'h4206e69c, 32'hc2c68703, 32'h4224aa15, 32'h41fe6cf5, 32'hc253d778, 32'hbf000586};
test_label[4381] = '{32'hc2c68703};
test_output[4381] = '{32'h430c7a21};
/*############ DEBUG ############
test_input[35048:35055] = '{38.1240226546, 29.1634880102, 33.7252046344, -99.2636970062, 41.1660966425, 31.8032007915, -52.9604185705, -0.500084257993};
test_label[4381] = '{-99.2636970062};
test_output[4381] = '{140.477072695};
############ END DEBUG ############*/
test_input[35056:35063] = '{32'hc29b6e7a, 32'h4289263f, 32'h4275ddb6, 32'h42402e86, 32'h40a561e9, 32'h40e0bdcd, 32'h42116d52, 32'h41e1eeaf};
test_label[4382] = '{32'h42402e86};
test_output[4382] = '{32'h41a43d9e};
/*############ DEBUG ############
test_input[35056:35063] = '{-77.7157737713, 68.5747026906, 61.4665146708, 48.045434951, 5.16820215689, 7.02316883258, 36.3567583961, 28.2415452718};
test_label[4382] = '{48.045434951};
test_output[4382] = '{20.5300857826};
############ END DEBUG ############*/
test_input[35064:35071] = '{32'hc2024911, 32'hc21c37c2, 32'h4175ec10, 32'h420d5e59, 32'hc1f2462f, 32'h40a784cf, 32'hc101ffbd, 32'hc20b8710};
test_label[4383] = '{32'h420d5e59};
test_output[4383] = '{32'h3111ab3e};
/*############ DEBUG ############
test_input[35064:35071] = '{-32.5713520573, -39.0544494042, 15.3701328854, 35.3421347255, -30.2842691675, 5.23496212184, -8.12493591591, -34.8818952213};
test_label[4383] = '{35.3421347255};
test_output[4383] = '{2.11976159073e-09};
############ END DEBUG ############*/
test_input[35072:35079] = '{32'hc299b826, 32'h42682763, 32'hc29a6043, 32'h42a0a25e, 32'hc23db1a6, 32'hc1e54c46, 32'h42bfb788, 32'h429160d3};
test_label[4384] = '{32'hc29a6043};
test_output[4384] = '{32'h432d0be6};
/*############ DEBUG ############
test_input[35072:35079] = '{-76.8596648865, 58.0384631882, -77.188011938, 80.3171236887, -47.4234849356, -28.6622438263, 95.8584619207, 72.6891062613};
test_label[4384] = '{-77.188011938};
test_output[4384] = '{173.046474037};
############ END DEBUG ############*/
test_input[35080:35087] = '{32'h42c7ce59, 32'h4235a408, 32'hc1ef80dc, 32'hc1a0d014, 32'h42187e6f, 32'h3f1d8dd8, 32'h42a07913, 32'hc2bfade1};
test_label[4385] = '{32'h42187e6f};
test_output[4385] = '{32'h42771e43};
/*############ DEBUG ############
test_input[35080:35087] = '{99.9030229862, 45.4101869769, -29.937918761, -20.1015999606, 38.1234697329, 0.615445616303, 80.2364722465, -95.8396106284};
test_label[4385] = '{38.1234697329};
test_output[4385] = '{61.7795532562};
############ END DEBUG ############*/
test_input[35088:35095] = '{32'hc1557efa, 32'hc2067028, 32'h42bdc514, 32'hc1800117, 32'h42b66ce8, 32'h41d2081b, 32'hc11d1722, 32'hc1bfc81a};
test_label[4386] = '{32'h41d2081b};
test_output[4386] = '{32'h42894fe7};
/*############ DEBUG ############
test_input[35088:35095] = '{-13.343500087, -33.6095270381, 94.884917184, -16.0005319114, 91.2127060817, 26.2539569728, -9.81814738724, -23.9727052549};
test_label[4386] = '{26.2539569728};
test_output[4386] = '{68.656062692};
############ END DEBUG ############*/
test_input[35096:35103] = '{32'hc0585d5a, 32'hc208bbd7, 32'hc29b76e8, 32'h40ad6816, 32'hc2c7d1a8, 32'h425c2d82, 32'h42800125, 32'hc20cc129};
test_label[4387] = '{32'hc0585d5a};
test_output[4387] = '{32'h4286c421};
/*############ DEBUG ############
test_input[35096:35103] = '{-3.38069773824, -34.1834390471, -77.7322375333, 5.41895569998, -99.9094879134, 55.0444402578, 64.0022344448, -35.1886318679};
test_label[4387] = '{-3.38069773824};
test_output[4387] = '{67.3830609046};
############ END DEBUG ############*/
test_input[35104:35111] = '{32'hc2a8fa65, 32'hc28c9c06, 32'h420e8ff8, 32'hc1a51493, 32'h4265d4b2, 32'h426b8d29, 32'hc228b9c4, 32'h42893888};
test_label[4388] = '{32'hc28c9c06};
test_output[4388] = '{32'h430aea4c};
/*############ DEBUG ############
test_input[35104:35111] = '{-84.4890487406, -70.304736033, 35.6405951186, -20.6350451817, 57.4577113041, 58.8878519429, -42.181413636, 68.6104096116};
test_label[4388] = '{-70.304736033};
test_output[4388] = '{138.915219895};
############ END DEBUG ############*/
test_input[35112:35119] = '{32'h40c8b7ad, 32'h42ab44a7, 32'hc27d82ef, 32'hc17922df, 32'hc24afdb2, 32'h40944da2, 32'hc1ca5bb5, 32'h41bfcd80};
test_label[4389] = '{32'h40c8b7ad};
test_output[4389] = '{32'h429eb92c};
/*############ DEBUG ############
test_input[35112:35119] = '{6.27242145558, 85.6340856808, -63.3778642849, -15.5710134388, -50.7477496979, 4.63447645744, -25.2947781003, 23.9753426997};
test_label[4389] = '{6.27242145558};
test_output[4389] = '{79.3616642252};
############ END DEBUG ############*/
test_input[35120:35127] = '{32'h429fc330, 32'hc2c19a20, 32'hc17dbe9e, 32'hc218e456, 32'hc2744490, 32'h420bf38f, 32'h4248bc6c, 32'h42164c32};
test_label[4390] = '{32'h429fc330};
test_output[4390] = '{32'h2a0ea000};
/*############ DEBUG ############
test_input[35120:35127] = '{79.8812285428, -96.8010255299, -15.8590374047, -38.2229859518, -61.0669548609, 34.9878496465, 50.1840075159, 37.5744103354};
test_label[4390] = '{79.8812285428};
test_output[4390] = '{1.2667644711e-13};
############ END DEBUG ############*/
test_input[35128:35135] = '{32'hc224eee9, 32'h410b471c, 32'hc2be124f, 32'h41f11bc7, 32'h41fffc32, 32'h428fa579, 32'h42bfdd99, 32'h3fc9663b};
test_label[4391] = '{32'h410b471c};
test_output[4391] = '{32'h42ae74b5};
/*############ DEBUG ############
test_input[35128:35135] = '{-41.2333115942, 8.70486079208, -95.0357552574, 30.13856344, 31.9981419656, 71.8231884739, 95.932807543, 1.57343237321};
test_label[4391] = '{8.70486079208};
test_output[4391] = '{87.227946751};
############ END DEBUG ############*/
test_input[35136:35143] = '{32'h41f06654, 32'h3d1fb659, 32'hc2656d32, 32'hc28747a8, 32'hc1d8552a, 32'h42b8d389, 32'h425d7622, 32'hc132828e};
test_label[4392] = '{32'h3d1fb659};
test_output[4392] = '{32'h42b8bf93};
/*############ DEBUG ############
test_input[35136:35143] = '{30.0499658411, 0.0389922600412, -57.3566346126, -67.6399545442, -27.0415831686, 92.4131570738, 55.3653623406, -11.1568738611};
test_label[4392] = '{0.0389922600412};
test_output[4392] = '{92.3741648137};
############ END DEBUG ############*/
test_input[35144:35151] = '{32'hc2538bec, 32'h3f5b3280, 32'h42c76fab, 32'h42bfd241, 32'h4269e3ff, 32'hc2accc77, 32'hbf8f7bc1, 32'hc2bb039c};
test_label[4393] = '{32'h3f5b3280};
test_output[4393] = '{32'h42c5c485};
/*############ DEBUG ############
test_input[35144:35151] = '{-52.8866411873, 0.856239343518, 99.7181029982, 95.9106522832, 58.4726513866, -86.3993429954, -1.12096413894, -93.5070505335};
test_label[4393] = '{0.856239343518};
test_output[4393] = '{98.8838254326};
############ END DEBUG ############*/
test_input[35152:35159] = '{32'hc1ea9ff3, 32'h42bc221a, 32'hc2a89d3a, 32'h41bd1c2f, 32'hc0e107d0, 32'h42bff7a8, 32'h429733e9, 32'hc2a78e26};
test_label[4394] = '{32'hc0e107d0};
test_output[4394] = '{32'h42ce4e62};
/*############ DEBUG ############
test_input[35152:35159] = '{-29.328099302, 94.0666067421, -84.3070797752, 23.6387609935, -7.03220348347, 95.9837060728, 75.6013876564, -83.7776374586};
test_label[4394] = '{-7.03220348347};
test_output[4394] = '{103.153088025};
############ END DEBUG ############*/
test_input[35160:35167] = '{32'hc2899de2, 32'hc2c72d31, 32'hc1deb87d, 32'hc1c844dd, 32'hc240c1c6, 32'hbe7e57f5, 32'hc27640bd, 32'h424fce3a};
test_label[4395] = '{32'hc2c72d31};
test_output[4395] = '{32'h43178a27};
/*############ DEBUG ############
test_input[35160:35167] = '{-68.8083645757, -99.588262896, -27.8400813943, -25.0336246472, -48.1892308859, -0.248382400905, -61.5632209583, 51.9513949007};
test_label[4395] = '{-99.588262896};
test_output[4395] = '{151.539657797};
############ END DEBUG ############*/
test_input[35168:35175] = '{32'h42046b3e, 32'h42bfd298, 32'h428cba6b, 32'hc16469c6, 32'hc215cf29, 32'hc2bb3f2e, 32'hc2647337, 32'hc2828203};
test_label[4396] = '{32'hc16469c6};
test_output[4396] = '{32'h42dc5fd1};
/*############ DEBUG ############
test_input[35168:35175] = '{33.1047298223, 95.911319192, 70.3640940871, -14.2758232312, -37.4523040794, -93.6234013533, -57.1125138948, -65.2539282372};
test_label[4396] = '{-14.2758232312};
test_output[4396] = '{110.187142423};
############ END DEBUG ############*/
test_input[35176:35183] = '{32'hc28aeb3d, 32'hc237413a, 32'h423b5605, 32'hc281ef04, 32'h41bde6b3, 32'hc1b646da, 32'hc2852511, 32'hc2c2d293};
test_label[4397] = '{32'hc2c2d293};
test_output[4397] = '{32'h43103ecb};
/*############ DEBUG ############
test_input[35176:35183] = '{-69.4594486039, -45.8136988693, 46.834004281, -64.9668241815, 23.7376464987, -22.7845961238, -66.5723944337, -97.4112770008};
test_label[4397] = '{-97.4112770008};
test_output[4397] = '{144.245281282};
############ END DEBUG ############*/
test_input[35184:35191] = '{32'hc2394900, 32'hc2715574, 32'h40aa3eeb, 32'hc2c6f5cd, 32'h42386e0b, 32'h428400db, 32'hc29fc9a9, 32'hbf9937b1};
test_label[4398] = '{32'hbf9937b1};
test_output[4398] = '{32'h428665b9};
/*############ DEBUG ############
test_input[35184:35191] = '{-46.3212886972, -60.3334503761, 5.32018037128, -99.480076021, 46.1074636688, 66.001668334, -79.8938641115, -1.19701209989};
test_label[4398] = '{-1.19701209989};
test_output[4398] = '{67.1986804362};
############ END DEBUG ############*/
test_input[35192:35199] = '{32'hc2c0f023, 32'h424aa234, 32'h41b4f591, 32'h428c748f, 32'hc2b109f1, 32'h4070ddda, 32'h42485fd4, 32'hc2292078};
test_label[4399] = '{32'h4070ddda};
test_output[4399] = '{32'h4284eda1};
/*############ DEBUG ############
test_input[35192:35199] = '{-96.4690180069, 50.6583998918, 22.619906076, 70.2276562245, -88.5194178274, 3.7635407585, 50.0935834202, -42.2817074242};
test_label[4399] = '{3.7635407585};
test_output[4399] = '{66.464115471};
############ END DEBUG ############*/
test_input[35200:35207] = '{32'hc294829d, 32'hc299c239, 32'h42af448a, 32'hc224f766, 32'h427809ab, 32'h4248e09c, 32'hc16a2649, 32'hc2766fa4};
test_label[4400] = '{32'hc224f766};
test_output[4400] = '{32'h4300e01f};
/*############ DEBUG ############
test_input[35200:35207] = '{-74.2551018787, -76.8793396766, 87.6338652034, -41.2416005756, 62.0094405398, 50.219343272, -14.6343465136, -61.6090237024};
test_label[4400] = '{-41.2416005756};
test_output[4400] = '{128.875465779};
############ END DEBUG ############*/
test_input[35208:35215] = '{32'h4129cef4, 32'h42b5f3ef, 32'h426ab17b, 32'h3fe53557, 32'h429ec3dd, 32'h429afd7a, 32'h40f6f818, 32'h42b76814};
test_label[4401] = '{32'h3fe53557};
test_output[4401] = '{32'h42b49d29};
/*############ DEBUG ############
test_input[35208:35215] = '{10.6130257066, 90.9764351324, 58.6733222621, 1.79069033402, 79.3825451688, 77.4950743595, 7.71778503128, 91.7032809928};
test_label[4401] = '{1.79069033402};
test_output[4401] = '{90.3069520357};
############ END DEBUG ############*/
test_input[35216:35223] = '{32'h42472b10, 32'h4129d54b, 32'h401c5945, 32'h42c00018, 32'h4218a2a9, 32'hc1f65780, 32'hc29fa264, 32'hc1b52e6a};
test_label[4402] = '{32'h42472b10};
test_output[4402] = '{32'h4238d520};
/*############ DEBUG ############
test_input[35216:35223] = '{49.7920548967, 10.6145737781, 2.44294852351, 96.0001842339, 38.1588486306, -30.792723742, -79.8171672151, -22.6476631225};
test_label[4402] = '{49.7920548967};
test_output[4402] = '{46.2081293372};
############ END DEBUG ############*/
test_input[35224:35231] = '{32'hc29acfe6, 32'h420a3979, 32'hc28fbe5b, 32'h4265e9c4, 32'hc194adbe, 32'h4136686e, 32'hc160382d, 32'h4222bcec};
test_label[4403] = '{32'h420a3979};
test_output[4403] = '{32'h41b76096};
/*############ DEBUG ############
test_input[35224:35231] = '{-77.4060505548, 34.5561269155, -71.8717904438, 57.4782878999, -18.5848349242, 11.4004956995, -14.0137144491, 40.6844936307};
test_label[4403] = '{34.5561269155};
test_output[4403] = '{22.9221610353};
############ END DEBUG ############*/
test_input[35232:35239] = '{32'h41c23dc6, 32'h42648aa1, 32'hc29cdf52, 32'hc1e56467, 32'h42b4bcbf, 32'h4292f003, 32'h41abb60c, 32'hc07ba43b};
test_label[4404] = '{32'hc1e56467};
test_output[4404] = '{32'h42ee15d8};
/*############ DEBUG ############
test_input[35232:35239] = '{24.2801628355, 57.1353799856, -78.4361707849, -28.6740251822, 90.3686410952, 73.4687698053, 21.4638893445, -3.93189884901};
test_label[4404] = '{-28.6740251822};
test_output[4404] = '{119.042666323};
############ END DEBUG ############*/
test_input[35240:35247] = '{32'h42c12177, 32'hc2c0e774, 32'hc22d3b3b, 32'h41ae94f5, 32'hc293c9fb, 32'hc23f1eac, 32'h419ae96f, 32'h42af627f};
test_label[4405] = '{32'hc2c0e774};
test_output[4405] = '{32'h4341047f};
/*############ DEBUG ############
test_input[35240:35247] = '{96.5653588307, -96.4520576555, -43.3078413316, 21.8227320116, -73.894493284, -47.779952128, 19.3639819467, 87.6923769375};
test_label[4405] = '{-96.4520576555};
test_output[4405] = '{193.017556601};
############ END DEBUG ############*/
test_input[35248:35255] = '{32'hc2b84f76, 32'hc19a196a, 32'hc249051f, 32'hc1857ff2, 32'h42b56614, 32'h40be9cdd, 32'hc26f0891, 32'h4195ea62};
test_label[4406] = '{32'hc26f0891};
test_output[4406] = '{32'h4316752e};
/*############ DEBUG ############
test_input[35248:35255] = '{-92.1551953709, -19.2624086572, -50.255000816, -16.6874736511, 90.6993678694, 5.95664846404, -59.7583668553, 18.7394441243};
test_label[4406] = '{-59.7583668553};
test_output[4406] = '{150.457734725};
############ END DEBUG ############*/
test_input[35256:35263] = '{32'h419b6e80, 32'hc1d13495, 32'hc2870d47, 32'hc2b1ec87, 32'hc272d00e, 32'hc08aaf12, 32'hc2494cd7, 32'hc26d7a8c};
test_label[4407] = '{32'hc08aaf12};
test_output[4407] = '{32'h41be1a45};
/*############ DEBUG ############
test_input[35256:35263] = '{19.4289559563, -26.1506751251, -67.5259291444, -88.9619664088, -60.7031767272, -4.33387095353, -50.3250393637, -59.3696753691};
test_label[4407] = '{-4.33387095353};
test_output[4407] = '{23.7628269099};
############ END DEBUG ############*/
test_input[35264:35271] = '{32'hc286d88b, 32'hc2809c7f, 32'hc29974a1, 32'hc1e9b5ab, 32'hc229b9e8, 32'hc2b84171, 32'hc2800e24, 32'h42b24d21};
test_label[4408] = '{32'hc229b9e8};
test_output[4408] = '{32'h4303950b};
/*############ DEBUG ############
test_input[35264:35271] = '{-67.4229383579, -64.3056598175, -76.727788504, -29.2137055111, -42.4315493492, -92.1278122932, -64.0276185504, 89.1506454213};
test_label[4408] = '{-42.4315493492};
test_output[4408] = '{131.58219477};
############ END DEBUG ############*/
test_input[35272:35279] = '{32'h41285ed0, 32'hc2c65402, 32'hc2b940c7, 32'hc281a370, 32'h4261b399, 32'hc1a33529, 32'hc2bddd51, 32'hc11181f7};
test_label[4409] = '{32'h4261b399};
test_output[4409] = '{32'h80000000};
/*############ DEBUG ############
test_input[35272:35279] = '{10.5231479314, -99.1640783425, -92.6265178363, -64.8192133304, 56.4253886488, -20.4009571497, -94.9322570064, -9.09422933682};
test_label[4409] = '{56.4253886488};
test_output[4409] = '{-0.0};
############ END DEBUG ############*/
test_input[35280:35287] = '{32'h3f74a250, 32'h427b8f50, 32'hc1514501, 32'h42bb7f0a, 32'hc23b3df6, 32'hc0831759, 32'h4207250a, 32'hc28af06c};
test_label[4410] = '{32'h427b8f50};
test_output[4410] = '{32'h41f6dd89};
/*############ DEBUG ############
test_input[35280:35287] = '{0.955601680095, 62.8899534162, -13.0793468531, 93.7481243233, -46.8105098804, -4.09659999429, 33.7861713538, -69.469575942};
test_label[4410] = '{62.8899534162};
test_output[4410] = '{30.8581709071};
############ END DEBUG ############*/
test_input[35288:35295] = '{32'hc23dcaca, 32'h42320135, 32'hc276c7d0, 32'hc2a551d6, 32'h4114cf64, 32'h42bf8e4a, 32'hc29b3a76, 32'hc09b596a};
test_label[4411] = '{32'hc09b596a};
test_output[4411] = '{32'h42c943e0};
/*############ DEBUG ############
test_input[35288:35295] = '{-47.448034787, 44.501179095, -61.6951288753, -82.6598393908, 9.30063217881, 95.7779068543, -77.6141841058, -4.85466500072};
test_label[4411] = '{-4.85466500072};
test_output[4411] = '{100.632571855};
############ END DEBUG ############*/
test_input[35296:35303] = '{32'h40c2eaa0, 32'h4205ccbc, 32'h41f23cba, 32'hbfd3b37a, 32'h422a9fd0, 32'h4260fc5b, 32'hc29ad937, 32'hc2463dd2};
test_label[4412] = '{32'h4260fc5b};
test_output[4412] = '{32'h35a81fe1};
/*############ DEBUG ############
test_input[35296:35303] = '{6.09114052022, 33.4499344111, 30.279652594, -1.65391466753, 42.656067329, 56.2464403123, -77.4242444197, -49.5603726947};
test_label[4412] = '{56.2464403123};
test_output[4412] = '{1.25262529066e-06};
############ END DEBUG ############*/
test_input[35304:35311] = '{32'hc2ae6f25, 32'hc213ca85, 32'hc0db4f31, 32'h42a615cc, 32'hc2c019bd, 32'h41fdd1f8, 32'h41e4ebf8, 32'h4258fb0c};
test_label[4413] = '{32'hc2c019bd};
test_output[4413] = '{32'h433317c4};
/*############ DEBUG ############
test_input[35304:35311] = '{-87.2170828262, -36.9477729972, -6.8534169064, 83.0425695674, -96.0502717998, 31.7275229026, 28.6152191113, 54.2451631469};
test_label[4413] = '{-96.0502717998};
test_output[4413] = '{179.092841367};
############ END DEBUG ############*/
test_input[35312:35319] = '{32'h41861544, 32'h422e628a, 32'h42bfde33, 32'hc1fa8085, 32'hc2b4f643, 32'hbf0ba4e7, 32'hc205487c, 32'h42af18be};
test_label[4414] = '{32'h41861544};
test_output[4414] = '{32'h429e5900};
/*############ DEBUG ############
test_input[35312:35319] = '{16.7603841711, 43.5962288601, 95.9339860744, -31.3127545142, -90.4809805964, -0.545484931935, -33.3207851432, 87.5483226162};
test_label[4414] = '{16.7603841711};
test_output[4414] = '{79.1738299917};
############ END DEBUG ############*/
test_input[35320:35327] = '{32'hc1118c53, 32'hc18ba5c6, 32'hc2aa6bd7, 32'hc20bb0f8, 32'hbf29c01f, 32'h42ad4dcd, 32'h4289f282, 32'h427b9a0c};
test_label[4415] = '{32'hc2aa6bd7};
test_output[4415] = '{32'h432bdcd2};
/*############ DEBUG ############
test_input[35320:35327] = '{-9.09675895557, -17.4559445269, -85.2106260133, -34.922819298, -0.663087796627, 86.6519517736, 68.9736463076, 62.9004372473};
test_label[4415] = '{-85.2106260133};
test_output[4415] = '{171.862577808};
############ END DEBUG ############*/
test_input[35328:35335] = '{32'h3febb0c2, 32'hc2c3d27a, 32'h4215a169, 32'hc2a4a889, 32'h42a1f528, 32'hc1a4bb54, 32'h4293291a, 32'hc2810295};
test_label[4416] = '{32'h4293291a};
test_output[4416] = '{32'h40ecc5e6};
/*############ DEBUG ############
test_input[35328:35335] = '{1.84133167489, -97.9110898737, 37.4076287845, -82.3291667, 80.9788239248, -20.591467997, 73.5802785362, -64.505040491};
test_label[4416] = '{73.5802785362};
test_output[4416] = '{7.3991573439};
############ END DEBUG ############*/
test_input[35336:35343] = '{32'h415fc831, 32'hc25cc818, 32'hc1b0ce17, 32'hc0352c61, 32'hc2a0c785, 32'h421d16b7, 32'hc29dd66a, 32'h4253b96f};
test_label[4417] = '{32'h415fc831};
test_output[4417] = '{32'h421bc763};
/*############ DEBUG ############
test_input[35336:35343] = '{13.9863749887, -55.1954050661, -22.1006304252, -2.83083356002, -80.3896900438, 39.2721821988, -78.9187743711, 52.931086225};
test_label[4417] = '{13.9863749887};
test_output[4417] = '{38.9447124058};
############ END DEBUG ############*/
test_input[35344:35351] = '{32'h424c9326, 32'h41ea037d, 32'hc15b6057, 32'hc29604a8, 32'h41ca87e2, 32'h42bc7007, 32'hc14c6287, 32'h426f3e14};
test_label[4418] = '{32'h424c9326};
test_output[4418] = '{32'h422c4ce8};
/*############ DEBUG ############
test_input[35344:35351] = '{51.1436998779, 29.2517025648, -13.7110201885, -75.0090910541, 25.3163488239, 94.2188047761, -12.7740548998, 59.8106232498};
test_label[4418] = '{51.1436998779};
test_output[4418] = '{43.0751048983};
############ END DEBUG ############*/
test_input[35352:35359] = '{32'hc294287f, 32'hc263404c, 32'hc143e452, 32'hc0516385, 32'h423c2e1a, 32'hc29431c6, 32'hbf62498c, 32'h420bc919};
test_label[4419] = '{32'h420bc919};
test_output[4419] = '{32'h4141940d};
/*############ DEBUG ############
test_input[35352:35359] = '{-74.0790923033, -56.8127891788, -12.2432421982, -3.27169920138, 47.0450223134, -74.09721308, -0.883934715715, 34.9463829106};
test_label[4419] = '{34.9463829106};
test_output[4419] = '{12.0986449699};
############ END DEBUG ############*/
test_input[35360:35367] = '{32'h42088d01, 32'h4100deb1, 32'h423a8890, 32'h42882052, 32'hc12e741b, 32'hc2871d32, 32'hc241182d, 32'h42b6e6eb};
test_label[4420] = '{32'h42b6e6eb};
test_output[4420] = '{32'h2e991b90};
/*############ DEBUG ############
test_input[35360:35367] = '{34.1377002301, 8.054368339, 46.6333599496, 68.0631226568, -10.9033464369, -67.5570213944, -48.2736088512, 91.4510145839};
test_label[4420] = '{91.4510145839};
test_output[4420] = '{6.96253055234e-11};
############ END DEBUG ############*/
test_input[35368:35375] = '{32'h42b0c886, 32'h426ed7b1, 32'h429f17ca, 32'hc23b7b3c, 32'hc227d6ce, 32'hc1ef434b, 32'h4259ea1d, 32'hc1c6097e};
test_label[4421] = '{32'hc23b7b3c};
test_output[4421] = '{32'h4307431c};
/*############ DEBUG ############
test_input[35368:35375] = '{88.391646969, 59.7106379535, 79.5464631397, -46.8703477255, -41.9597683484, -29.9078571867, 54.4786247883, -24.7546343948};
test_label[4421] = '{-46.8703477255};
test_output[4421] = '{135.262138758};
############ END DEBUG ############*/
test_input[35376:35383] = '{32'h428beebd, 32'h41fec547, 32'hc19d66ff, 32'h408101af, 32'hc2b58689, 32'h42a65eea, 32'h427de9c0, 32'hc25ea16f};
test_label[4422] = '{32'hc25ea16f};
test_output[4422] = '{32'h430ad7d1};
/*############ DEBUG ############
test_input[35376:35383] = '{69.9662850053, 31.8463270048, -19.6752907023, 4.03145534024, -90.7627611064, 83.185381724, 63.4782718702, -55.657651441};
test_label[4422] = '{-55.657651441};
test_output[4422] = '{138.843034983};
############ END DEBUG ############*/
test_input[35384:35391] = '{32'hc1a7bf3a, 32'hc2b89100, 32'hc2bc7119, 32'hc29d06f9, 32'hc26716b9, 32'h42c3f256, 32'hc18913ad, 32'h4296553c};
test_label[4423] = '{32'hc2bc7119};
test_output[4423] = '{32'h434031b7};
/*############ DEBUG ############
test_input[35384:35391] = '{-20.9683718242, -92.2832028834, -94.2208930485, -78.5136166729, -57.7721916106, 97.973310083, -17.1346063762, 75.1664744793};
test_label[4423] = '{-94.2208930485};
test_output[4423] = '{192.194203132};
############ END DEBUG ############*/
test_input[35392:35399] = '{32'h425a6fd0, 32'h42a61c3c, 32'h41b58c20, 32'hc09a5fa0, 32'h423ad3f7, 32'h40af70fb, 32'h40123de7, 32'hc2c408a5};
test_label[4424] = '{32'h41b58c20};
test_output[4424] = '{32'h42717269};
/*############ DEBUG ############
test_input[35392:35399] = '{54.6091923101, 83.0551477415, 22.6934205067, -4.82417287677, 46.7069972979, 5.48254133058, 2.28502826785, -98.0168858121};
test_label[4424] = '{22.6934205067};
test_output[4424] = '{60.3617272348};
############ END DEBUG ############*/
test_input[35400:35407] = '{32'hc2ac37d3, 32'hc2aa2be1, 32'h428abeb5, 32'hc2484ae5, 32'h42c7bc35, 32'h418236e0, 32'hc17f5e9d, 32'hc22802f6};
test_label[4425] = '{32'hc17f5e9d};
test_output[4425] = '{32'h42e7a809};
/*############ DEBUG ############
test_input[35400:35407] = '{-86.1090316346, -85.0856995732, 69.3724773849, -50.0731392567, 99.8675916349, 16.2767952346, -15.9605986547, -42.0028932167};
test_label[4425] = '{-15.9605986547};
test_output[4425] = '{115.82819029};
############ END DEBUG ############*/
test_input[35408:35415] = '{32'hc27f55a4, 32'hc29ebaf9, 32'hc1abe4c3, 32'hc296d3c2, 32'h428f5a5c, 32'h4209da32, 32'h41fc69ba, 32'h41606545};
test_label[4426] = '{32'hc27f55a4};
test_output[4426] = '{32'h43078297};
/*############ DEBUG ############
test_input[35408:35415] = '{-63.83363385, -79.3651843825, -21.4866998879, -75.4135912831, 71.676482653, 34.4630823223, 31.5516249446, 14.0247236467};
test_label[4426] = '{-63.83363385};
test_output[4426] = '{135.510116503};
############ END DEBUG ############*/
test_input[35416:35423] = '{32'h429e2dcc, 32'hc1ff3238, 32'hc2643157, 32'hc19db9ab, 32'h4259c26d, 32'h41504e20, 32'h42b3b059, 32'hc16c0dd6};
test_label[4427] = '{32'h41504e20};
test_output[4427] = '{32'h4299a698};
/*############ DEBUG ############
test_input[35416:35423] = '{79.0894494179, -31.8995210199, -57.0481841813, -19.7156574296, 54.4398697585, 13.0190738686, 89.8444282843, -14.7533781797};
test_label[4427] = '{13.0190738686};
test_output[4427] = '{76.8253757544};
############ END DEBUG ############*/
test_input[35424:35431] = '{32'hc08a3c78, 32'hc2b0893f, 32'h41f148c5, 32'h41009e39, 32'h42aed318, 32'h4216abe6, 32'h42a4441e, 32'hbec03692};
test_label[4428] = '{32'h42aed318};
test_output[4428] = '{32'h3ba691f3};
/*############ DEBUG ############
test_input[35424:35431] = '{-4.31988126789, -88.2680595161, 30.1605325811, 8.03862816119, 87.4122936271, 37.6678687128, 82.1330449743, -0.375416336808};
test_label[4428] = '{87.4122936271};
test_output[4428] = '{0.00508331644092};
############ END DEBUG ############*/
test_input[35432:35439] = '{32'h42a88a3a, 32'hc1a9db10, 32'h408415a6, 32'hc27a820b, 32'hc24b9417, 32'h422f8be6, 32'h42a1fafe, 32'hc28b8619};
test_label[4429] = '{32'hc1a9db10};
test_output[4429] = '{32'h42d313e9};
/*############ DEBUG ############
test_input[35432:35439] = '{84.2699772896, -21.2319635329, 4.12764263314, -62.6269941698, -50.8946205372, 43.8866187795, 80.9902178948, -69.7619088641};
test_label[4429] = '{-21.2319635329};
test_output[4429] = '{105.538887135};
############ END DEBUG ############*/
test_input[35440:35447] = '{32'h419eb166, 32'h4253fb01, 32'hbfba0fef, 32'h425942c8, 32'hc209390a, 32'h41aaf497, 32'h42a77f4a, 32'h421a13f1};
test_label[4430] = '{32'h419eb166};
test_output[4430] = '{32'h427fa5e1};
/*############ DEBUG ############
test_input[35440:35447] = '{19.836619698, 52.9951197998, -1.45361122008, 54.3152171034, -34.305703363, 21.3694286883, 83.7486096597, 38.5194749483};
test_label[4430] = '{19.836619698};
test_output[4430] = '{63.9119899617};
############ END DEBUG ############*/
test_input[35448:35455] = '{32'hc2b6e2c8, 32'hc297cae5, 32'h41f092ee, 32'hc16c28b7, 32'hc2928199, 32'hc188dd0f, 32'h4250431a, 32'hc1c339ea};
test_label[4431] = '{32'hc16c28b7};
test_output[4431] = '{32'h4285a6a4};
/*############ DEBUG ############
test_input[35448:35455] = '{-91.4429326748, -75.8962763057, 30.0717424265, -14.7599404311, -73.2531205825, -17.107937878, 52.0655298351, -24.4032788669};
test_label[4431] = '{-14.7599404311};
test_output[4431] = '{66.8254702665};
############ END DEBUG ############*/
test_input[35456:35463] = '{32'h405ce578, 32'h41b658bf, 32'h427db24b, 32'hc2c547ea, 32'hc1a643c8, 32'hc0befe60, 32'h42b1f21f, 32'h42a22194};
test_label[4432] = '{32'h42a22194};
test_output[4432] = '{32'h40fd0bae};
/*############ DEBUG ############
test_input[35456:35463] = '{3.45150565729, 22.793332783, 63.4241147099, -98.6404535912, -20.7830971687, -5.9685514146, 88.9728910836, 81.0655830838};
test_label[4432] = '{81.0655830838};
test_output[4432] = '{7.9076759762};
############ END DEBUG ############*/
test_input[35464:35471] = '{32'hc2b668ea, 32'h42babaa0, 32'hc2189159, 32'h41e4f2e9, 32'hc2122bd0, 32'hc2aaf2bd, 32'h419e1ace, 32'h42561300};
test_label[4433] = '{32'hc2aaf2bd};
test_output[4433] = '{32'h4332d6ae};
/*############ DEBUG ############
test_input[35464:35471] = '{-91.2049093277, 93.3645011931, -38.1419392632, 28.618608239, -36.5427841708, -85.4740952279, 19.7630888766, 53.5185559553};
test_label[4433] = '{-85.4740952279};
test_output[4433] = '{178.838596421};
############ END DEBUG ############*/
test_input[35472:35479] = '{32'hc21d6a77, 32'h42b9e3f3, 32'hc1d533fb, 32'hc25d4414, 32'hc21523e3, 32'h41c75746, 32'hc1f7303a, 32'hc252f90e};
test_label[4434] = '{32'hc1d533fb};
test_output[4434] = '{32'h42ef30f2};
/*############ DEBUG ############
test_input[35472:35479] = '{-39.3539698381, 92.9452150984, -26.6503816507, -55.3164816834, -37.285047346, 24.9176138009, -30.8985486263, -52.7432184806};
test_label[4434] = '{-26.6503816507};
test_output[4434] = '{119.595596749};
############ END DEBUG ############*/
test_input[35480:35487] = '{32'h42ab8752, 32'h41748c31, 32'h42bf2ffa, 32'hc1bbee0c, 32'h42b6a057, 32'h42358722, 32'h42b2f5aa, 32'hc1c8bc61};
test_label[4435] = '{32'h42bf2ffa};
test_output[4435] = '{32'h3c82d957};
/*############ DEBUG ############
test_input[35480:35487] = '{85.7642950927, 15.2842261394, 95.5937031179, -23.4912344048, 91.3131674982, 45.3819666966, 89.4798125766, -25.0919812329};
test_label[4435] = '{95.5937031179};
test_output[4435] = '{0.0159727760483};
############ END DEBUG ############*/
test_input[35488:35495] = '{32'hc29fee2f, 32'h42acac93, 32'hbf11cf9c, 32'hc12aeb0f, 32'h427a1d5d, 32'h42b0557c, 32'h42b1e7f7, 32'hc297a0b2};
test_label[4436] = '{32'hc297a0b2};
test_output[4436] = '{32'h432530fc};
/*############ DEBUG ############
test_input[35488:35495] = '{-79.9651990554, 86.3370621167, -0.569574089635, -10.6823876611, 62.5286743177, 88.1669626709, 88.9530545203, -75.8138564257};
test_label[4436] = '{-75.8138564257};
test_output[4436] = '{165.19133988};
############ END DEBUG ############*/
test_input[35496:35503] = '{32'hc226c795, 32'h423787ba, 32'hc2b553a8, 32'hc261e52d, 32'hc2b8f84d, 32'h42a54a74, 32'h3f2e8e54, 32'h422ba3f5};
test_label[4437] = '{32'h3f2e8e54};
test_output[4437] = '{32'h42a3ed57};
/*############ DEBUG ############
test_input[35496:35503] = '{-41.6949060394, 45.8825437348, -90.663388366, -56.473804938, -92.4849657252, 82.6454136655, 0.681859237631, 42.9101152531};
test_label[4437] = '{0.681859237631};
test_output[4437] = '{81.9635544279};
############ END DEBUG ############*/
test_input[35504:35511] = '{32'hc21213e7, 32'hc2bef576, 32'hc24579ef, 32'h4265a25b, 32'h42810ede, 32'h42311324, 32'h41845790, 32'h4286fa8f};
test_label[4438] = '{32'h4286fa8f};
test_output[4438] = '{32'h3d4f0738};
/*############ DEBUG ############
test_input[35504:35511] = '{-36.5194371711, -95.4794152422, -49.3690743044, 57.4085499474, 64.5290348009, 44.2686920036, 16.5427545397, 67.4893755816};
test_label[4438] = '{67.4893755816};
test_output[4438] = '{0.0505439931279};
############ END DEBUG ############*/
test_input[35512:35519] = '{32'hc28fef19, 32'hc2847765, 32'h41ae34cc, 32'hc20b1cde, 32'h41532f32, 32'hc1c805e9, 32'hc299c32e, 32'h42111ab1};
test_label[4439] = '{32'hc1c805e9};
test_output[4439] = '{32'h42751da6};
/*############ DEBUG ############
test_input[35512:35519] = '{-71.9669858166, -66.2331952633, 21.7757794777, -34.7781892052, 13.199021974, -25.0028859129, -76.8812082877, 36.2760664327};
test_label[4439] = '{-25.0028859129};
test_output[4439] = '{61.2789528499};
############ END DEBUG ############*/
test_input[35520:35527] = '{32'hc2bc5f15, 32'hc08484a2, 32'h41d7f62b, 32'hc0e3c7b4, 32'h4281dbf0, 32'h4242af6a, 32'h4232765e, 32'hc12ddcc3};
test_label[4440] = '{32'hc12ddcc3};
test_output[4440] = '{32'h42979788};
/*############ DEBUG ############
test_input[35520:35527] = '{-94.1857048493, -4.14119033126, 26.9952000735, -7.11812758646, 64.9295643386, 48.6713020327, 44.6155939692, -10.86639704};
test_label[4440] = '{-10.86639704};
test_output[4440] = '{75.7959614671};
############ END DEBUG ############*/
test_input[35528:35535] = '{32'h425015f0, 32'h41d4fbb5, 32'hc2bd18ae, 32'h4287b75b, 32'h42c44f9f, 32'hc23cb037, 32'hc196eb9a, 32'hc2380a10};
test_label[4441] = '{32'h4287b75b};
test_output[4441] = '{32'h41f26110};
/*############ DEBUG ############
test_input[35528:35535] = '{52.0214224348, 26.6229034901, -94.54820136, 67.8581179351, 98.1555121767, -47.1720832651, -18.8650391411, -46.0098275725};
test_label[4441] = '{67.8581179351};
test_output[4441] = '{30.2973942415};
############ END DEBUG ############*/
test_input[35536:35543] = '{32'hc23ee72a, 32'hc23ef5ea, 32'hc0a910a7, 32'hc29d5f83, 32'h41d09a08, 32'h4163c03e, 32'h42819876, 32'h418af179};
test_label[4442] = '{32'h41d09a08};
test_output[4442] = '{32'h421ae3e8};
/*############ DEBUG ############
test_input[35536:35543] = '{-47.7257468385, -47.7401502189, -5.28328282142, -78.6865487339, 26.0752102257, 14.2344340226, 64.7977757869, 17.3679056742};
test_label[4442] = '{26.0752102257};
test_output[4442] = '{38.7225655611};
############ END DEBUG ############*/
test_input[35544:35551] = '{32'h418bd5fb, 32'hc2960c0a, 32'h427a004b, 32'hc29b988b, 32'h42bd82c1, 32'hc2c2e599, 32'hc191bc98, 32'h424733e5};
test_label[4443] = '{32'hc29b988b};
test_output[4443] = '{32'h432c8da6};
/*############ DEBUG ############
test_input[35544:35551] = '{17.4794822547, -75.0235120747, 62.5002844336, -77.7979389948, 94.7553784528, -97.4484333135, -18.2170869389, 49.8006777981};
test_label[4443] = '{-77.7979389948};
test_output[4443] = '{172.553317448};
############ END DEBUG ############*/
test_input[35552:35559] = '{32'hc2064750, 32'h41075bd2, 32'h4251f66a, 32'hc2c7babc, 32'hc0500e12, 32'hc234319c, 32'hc20d78e4, 32'hc297574d};
test_label[4444] = '{32'hc20d78e4};
test_output[4444] = '{32'h42afb7a7};
/*############ DEBUG ############
test_input[35552:35559] = '{-33.5696422645, 8.45991669607, 52.4906378102, -99.8647171319, -3.25085876106, -45.0484485076, -35.3680576904, -75.6705099827};
test_label[4444] = '{-35.3680576904};
test_output[4444] = '{87.8586955006};
############ END DEBUG ############*/
test_input[35560:35567] = '{32'h426705ea, 32'hc251ef8d, 32'hc0db796d, 32'h424c426d, 32'hc2a16dd4, 32'hc2b998de, 32'hc291bd46, 32'h429856d8};
test_label[4445] = '{32'hc2a16dd4};
test_output[4445] = '{32'h431ce256};
/*############ DEBUG ############
test_input[35560:35567] = '{57.7557746058, -52.4839369664, -6.85857239748, 51.0648672344, -80.7145067529, -92.7985719108, -72.8696745682, 76.1696169736};
test_label[4445] = '{-80.7145067529};
test_output[4445] = '{156.884123737};
############ END DEBUG ############*/
test_input[35568:35575] = '{32'hc0b4540d, 32'hc1a9b5e2, 32'h41f10fe6, 32'h4271473f, 32'hc29bd0b4, 32'h4257b1b2, 32'hc2817110, 32'h424de9dd};
test_label[4446] = '{32'hc2817110};
test_output[4446] = '{32'h42fa159c};
/*############ DEBUG ############
test_input[35568:35575] = '{-5.63526003421, -21.2138100615, 30.1327623489, 60.3195747791, -77.9076237582, 53.9235322092, -64.7208228209, 51.4783820018};
test_label[4446] = '{-64.7208228209};
test_output[4446] = '{125.042208755};
############ END DEBUG ############*/
test_input[35576:35583] = '{32'hc09bb1bf, 32'h41c871ab, 32'hc20907f5, 32'h429d90cc, 32'hc1ac5508, 32'hc1d5073e, 32'hc2489119, 32'hc2be3183};
test_label[4447] = '{32'hc2be3183};
test_output[4447] = '{32'h432de128};
/*############ DEBUG ############
test_input[35576:35583] = '{-4.86544768088, 25.0555010237, -34.2577724309, 78.782807493, -21.5415184106, -26.6285371506, -50.1416952732, -95.0967017435};
test_label[4447] = '{-95.0967017435};
test_output[4447] = '{173.879509237};
############ END DEBUG ############*/
test_input[35584:35591] = '{32'hc2267fc8, 32'hc25157f5, 32'hc2584cad, 32'h4282155c, 32'hc2948b79, 32'hc275ecef, 32'h426d8ce5, 32'hc1e5eb6e};
test_label[4448] = '{32'hc2267fc8};
test_output[4448] = '{32'h42d5570b};
/*############ DEBUG ############
test_input[35584:35591] = '{-41.6247862534, -52.3358955631, -54.074878639, 65.0417212189, -74.2724073612, -61.4813822365, 59.3875918366, -28.7399559302};
test_label[4448] = '{-41.6247862534};
test_output[4448] = '{106.670004373};
############ END DEBUG ############*/
test_input[35592:35599] = '{32'hc2582944, 32'h4280f73b, 32'hc0d5e1b8, 32'h4174f784, 32'hc1c51dc9, 32'hc203b64b, 32'hc26bb1de, 32'hc2798373};
test_label[4449] = '{32'hc0d5e1b8};
test_output[4449] = '{32'h428e5556};
/*############ DEBUG ############
test_input[35592:35599] = '{-54.0402990031, 64.4828689483, -6.68380361922, 15.3104290645, -24.6395430422, -32.9280201345, -58.9236982709, -62.3783690615};
test_label[4449] = '{-6.68380361922};
test_output[4449] = '{71.1666725675};
############ END DEBUG ############*/
test_input[35600:35607] = '{32'h423355c0, 32'h428b9d66, 32'hc0c05368, 32'h4214dbc6, 32'hc2aa422b, 32'h42269e83, 32'hc29b0a79, 32'h42654038};
test_label[4450] = '{32'h423355c0};
test_output[4450] = '{32'h41c7ca1a};
/*############ DEBUG ############
test_input[35600:35607] = '{44.8337412022, 69.807420333, -6.0101815287, 37.2146228624, -85.1292319835, 41.6547974568, -77.5204563225, 57.3127137114};
test_label[4450] = '{44.8337412022};
test_output[4450] = '{24.9736828773};
############ END DEBUG ############*/
test_input[35608:35615] = '{32'hc29ca7b5, 32'h410d9065, 32'hc1201e71, 32'hc1aa4a97, 32'hc2ab6655, 32'hc2471eab, 32'hc1fcee13, 32'hc2c17a3d};
test_label[4451] = '{32'hc2c17a3d};
test_output[4451] = '{32'h42d32c4a};
/*############ DEBUG ############
test_input[35608:35615] = '{-78.3275522136, 8.84775259352, -10.0074320263, -21.2864204052, -85.6998670882, -49.7799493082, -31.6162464385, -96.7387495722};
test_label[4451] = '{-96.7387495722};
test_output[4451] = '{105.586502172};
############ END DEBUG ############*/
test_input[35616:35623] = '{32'h40983396, 32'h42109c3d, 32'hc2b88fab, 32'h428a982b, 32'hc28e3bb9, 32'hc05ad928, 32'hbf06e8eb, 32'h429dfc5b};
test_label[4452] = '{32'h428a982b};
test_output[4452] = '{32'h411b21bd};
/*############ DEBUG ############
test_input[35616:35623] = '{4.75629721054, 36.1525772621, -92.2806005406, 69.2972034651, -71.1166427053, -3.41950413838, -0.526991573725, 78.9928788399};
test_label[4452] = '{69.2972034651};
test_output[4452] = '{9.69573692199};
############ END DEBUG ############*/
test_input[35624:35631] = '{32'hc266a9e3, 32'hc2ba5d7e, 32'h42c23d31, 32'h42a06d46, 32'hc2ae5322, 32'hc1d575fc, 32'hc22a7c1f, 32'h429f2785};
test_label[4453] = '{32'h42c23d31};
test_output[4453] = '{32'h339558be};
/*############ DEBUG ############
test_input[35624:35631] = '{-57.6659056315, -93.1825984172, 97.119514436, 80.2134257886, -87.1623691084, -26.682608936, -42.6212110183, 79.5771855647};
test_label[4453] = '{97.119514436};
test_output[4453] = '{6.95449505519e-08};
############ END DEBUG ############*/
test_input[35632:35639] = '{32'h42c2204b, 32'h42a2086c, 32'h42aafdb1, 32'hc24aa696, 32'hc10bb624, 32'h4293b0ed, 32'hc2892d21, 32'hc2be1757};
test_label[4454] = '{32'hc10bb624};
test_output[4454] = '{32'h42d39711};
/*############ DEBUG ############
test_input[35632:35639] = '{97.0630730549, 81.0164459311, 85.4954944403, -50.6626819614, -8.73196833759, 73.8455605452, -68.5881444361, -95.0455825828};
test_label[4454] = '{-8.73196833759};
test_output[4454] = '{105.795050968};
############ END DEBUG ############*/
test_input[35640:35647] = '{32'hc23413e3, 32'h41ec06cc, 32'h42a69d69, 32'hc1687cb6, 32'hc2ae9f91, 32'hc210461f, 32'hc2bb5d32, 32'hc2648d5d};
test_label[4455] = '{32'h41ec06cc};
test_output[4455] = '{32'h4257376c};
/*############ DEBUG ############
test_input[35640:35647] = '{-45.0194215989, 29.5033181995, 83.3074414346, -14.5304473225, -87.3116540295, -36.0684785505, -93.6820217025, -57.1380511563};
test_label[4455] = '{29.5033181995};
test_output[4455] = '{53.804123235};
############ END DEBUG ############*/
test_input[35648:35655] = '{32'hc152d5ba, 32'hc2a967ae, 32'h418f2aae, 32'h42994a36, 32'h42b97173, 32'hc2758d55, 32'hc16970c8, 32'h42747fe7};
test_label[4456] = '{32'h42994a36};
test_output[4456] = '{32'h41809cf4};
/*############ DEBUG ############
test_input[35648:35655] = '{-13.1771796274, -84.7024963144, 17.895839795, 76.6449446929, 92.7215812692, -61.3880208574, -14.5900341154, 61.124906418};
test_label[4456] = '{76.6449446929};
test_output[4456] = '{16.0766366805};
############ END DEBUG ############*/
test_input[35656:35663] = '{32'h425e032a, 32'hc1d4c5a7, 32'h42827d26, 32'hc28188b4, 32'hc25491a3, 32'h42471f26, 32'hc1582382, 32'h426321f5};
test_label[4457] = '{32'h425e032a};
test_output[4457] = '{32'h411bdda6};
/*############ DEBUG ############
test_input[35656:35663] = '{55.5030890159, -26.596509195, 65.2444317079, -64.7669997793, -53.1422222031, 49.7804189659, -13.5086690744, 56.783159341};
test_label[4457] = '{55.5030890159};
test_output[4457] = '{9.74161315214};
############ END DEBUG ############*/
test_input[35664:35671] = '{32'hc2343284, 32'hc185ab4c, 32'hc2b9b02b, 32'h3ecc5ee4, 32'h419fab75, 32'hc29e434c, 32'h42c18244, 32'h42bbcef2};
test_label[4458] = '{32'h42c18244};
test_output[4458] = '{32'h3d66479d};
/*############ DEBUG ############
test_input[35664:35671] = '{-45.0493322611, -16.708640325, -92.8440784871, 0.399161450907, 19.9587191976, -79.1314408589, 96.7544217756, 93.9041924653};
test_label[4458] = '{96.7544217756};
test_output[4458] = '{0.0562206402473};
############ END DEBUG ############*/
test_input[35672:35679] = '{32'h42ae809f, 32'h420888d6, 32'hc18bca89, 32'hc19428df, 32'hc2ad093a, 32'hc29d48b7, 32'hc275bf86, 32'hc25be1e8};
test_label[4459] = '{32'hc29d48b7};
test_output[4459] = '{32'h4325e4ab};
/*############ DEBUG ############
test_input[35672:35679] = '{87.2512094936, 34.1336273962, -17.4738946149, -18.5199558161, -86.5180168568, -78.642023296, -61.43703432, -54.9706131979};
test_label[4459] = '{-78.642023296};
test_output[4459] = '{165.89323279};
############ END DEBUG ############*/
test_input[35680:35687] = '{32'h42b4606c, 32'h42c0ee32, 32'h4209dd3f, 32'hc2acc4ba, 32'h42c1d209, 32'hc1f87c04, 32'hc20ccfd5, 32'hc18c2349};
test_label[4460] = '{32'hc2acc4ba};
test_output[4460] = '{32'h4337ca57};
/*############ DEBUG ############
test_input[35680:35687] = '{90.1883219114, 96.4652253342, 34.4660615421, -86.3842334543, 96.9102252711, -31.0605547816, -35.2029592232, -17.5172281826};
test_label[4460] = '{-86.3842334543};
test_output[4460] = '{183.79039113};
############ END DEBUG ############*/
test_input[35688:35695] = '{32'hbe1b11ed, 32'hc221d373, 32'hc17c9e1e, 32'h41746f9a, 32'hc2b04001, 32'h427f8d8a, 32'h424313f5, 32'hc28679f3};
test_label[4461] = '{32'hc17c9e1e};
test_output[4461] = '{32'h429f5a89};
/*############ DEBUG ############
test_input[35688:35695] = '{-0.151435563149, -40.4564924525, -15.7886025409, 15.2772463345, -88.1250096679, 63.8882214574, 48.7694892006, -67.2381813311};
test_label[4461] = '{-15.7886025409};
test_output[4461] = '{79.67682427};
############ END DEBUG ############*/
test_input[35696:35703] = '{32'hc2a6f814, 32'hc050b816, 32'h427e3ff8, 32'hc2a8b8ed, 32'hc2430272, 32'hc107b27f, 32'h42c6429e, 32'hc20bbb68};
test_label[4462] = '{32'h42c6429e};
test_output[4462] = '{32'h26000000};
/*############ DEBUG ############
test_input[35696:35703] = '{-83.4845243717, -3.26123570061, 63.5624690882, -84.3611797731, -48.7523889245, -8.48107794621, 99.130108876, -34.9330145874};
test_label[4462] = '{99.130108876};
test_output[4462] = '{4.4408920985e-16};
############ END DEBUG ############*/
test_input[35704:35711] = '{32'hc2ac9d3e, 32'h426afa80, 32'hc18c6bfe, 32'h41b00a0b, 32'h41a12f27, 32'h42ad9969, 32'h41e1970a, 32'h41b84f93};
test_label[4463] = '{32'hc18c6bfe};
test_output[4463] = '{32'h42d0b468};
/*############ DEBUG ############
test_input[35704:35711] = '{-86.30711078, 58.7446292412, -17.5527300813, 22.0049037164, 20.1480244813, 86.799627684, 28.1987503342, 23.0388549078};
test_label[4463] = '{-17.5527300813};
test_output[4463] = '{104.352357765};
############ END DEBUG ############*/
test_input[35712:35719] = '{32'hc158681c, 32'hc28e17a3, 32'hc23092c3, 32'hc1d4b667, 32'h411d42a0, 32'hc28b2ebf, 32'h41029270, 32'hc20317d3};
test_label[4464] = '{32'hc23092c3};
test_output[4464] = '{32'h4258945c};
/*############ DEBUG ############
test_input[35712:35719] = '{-13.5254171628, -71.0461662807, -44.1433235333, -26.5890639053, 9.82876609721, -69.5913036619, 8.16075159718, -32.7732656664};
test_label[4464] = '{-44.1433235333};
test_output[4464] = '{54.1448836117};
############ END DEBUG ############*/
test_input[35720:35727] = '{32'hc212f88b, 32'hc0a0b4e6, 32'h4140e997, 32'hc24ae89e, 32'h42b41245, 32'hc22753e8, 32'hc2a549b7, 32'hc282761c};
test_label[4465] = '{32'h4140e997};
test_output[4465] = '{32'h429bf512};
/*############ DEBUG ############
test_input[35720:35727] = '{-36.7427163449, -5.02208242215, 12.0570287958, -50.7271669297, 90.0356846101, -41.8319392802, -82.6439768682, -65.2306843737};
test_label[4465] = '{12.0570287958};
test_output[4465] = '{77.9786558144};
############ END DEBUG ############*/
test_input[35728:35735] = '{32'h41c7fb1b, 32'h428e3b7f, 32'hc27ee7f1, 32'h428b8efd, 32'h41571b1b, 32'hc22f835f, 32'h4268483a, 32'h4259ae35};
test_label[4466] = '{32'h428e3b7f};
test_output[4466] = '{32'h3e6ed024};
/*############ DEBUG ############
test_input[35728:35735] = '{24.9976102081, 71.1162029298, -63.7265049255, 69.7792768264, 13.4441178203, -43.8782930952, 58.0705330671, 54.4201236996};
test_label[4466] = '{71.1162029298};
test_output[4466] = '{0.233215862028};
############ END DEBUG ############*/
test_input[35736:35743] = '{32'hc28147b2, 32'hc207d559, 32'hc27e1243, 32'hc23837ce, 32'h419570a6, 32'hc1f060ab, 32'hc260689b, 32'hc2773f32};
test_label[4467] = '{32'h419570a6};
test_output[4467] = '{32'h80000000};
/*############ DEBUG ############
test_input[35736:35743] = '{-64.6400328358, -33.9583489593, -63.5178324316, -46.0544961912, 18.6800047402, -30.0472008844, -56.1021528534, -61.8117128107};
test_label[4467] = '{18.6800047402};
test_output[4467] = '{-0.0};
############ END DEBUG ############*/
test_input[35744:35751] = '{32'hc2c1f2bb, 32'h42a779d7, 32'hc1c58f61, 32'hc0e40c90, 32'hc2117a48, 32'h41ffdb90, 32'h4294a2fa, 32'hc28dbafc};
test_label[4468] = '{32'h4294a2fa};
test_output[4468] = '{32'h4116b73d};
/*############ DEBUG ############
test_input[35744:35751] = '{-96.9740820214, 83.7379667363, -24.6950101219, -7.12653347471, -36.3694159235, 31.9822081843, 74.3183117321, -70.8652054472};
test_label[4468] = '{74.3183117321};
test_output[4468] = '{9.41973611492};
############ END DEBUG ############*/
test_input[35752:35759] = '{32'hc240d746, 32'h42bdeed1, 32'hc19a5643, 32'hc204211a, 32'hc24f86c0, 32'hc1cda963, 32'h42488f5b, 32'hc297e128};
test_label[4469] = '{32'hc1cda963};
test_output[4469] = '{32'h42f1592a};
/*############ DEBUG ############
test_input[35752:35759] = '{-48.210226923, 94.9664379475, -19.2921190575, -33.0323270231, -51.8815926889, -25.7077074176, 50.1399949915, -75.9397578123};
test_label[4469] = '{-25.7077074176};
test_output[4469] = '{120.674145365};
############ END DEBUG ############*/
test_input[35760:35767] = '{32'hc2542830, 32'hc203418e, 32'hc248ec18, 32'h409e4523, 32'hc2b7b86a, 32'h425b97dc, 32'hc299236f, 32'hc23b824a};
test_label[4470] = '{32'hc23b824a};
test_output[4470] = '{32'h42cb8d13};
/*############ DEBUG ############
test_input[35760:35767] = '{-53.0392458941, -32.814017334, -50.2305607584, 4.94593933248, -91.8601831879, 54.898301381, -76.5692096104, -46.8772355787};
test_label[4470] = '{-46.8772355787};
test_output[4470] = '{101.77553696};
############ END DEBUG ############*/
test_input[35768:35775] = '{32'h3f8afa97, 32'h42b75b84, 32'h41aef84d, 32'h41357bc5, 32'h4079a63d, 32'hc230068c, 32'hc06423a7, 32'h4182d38a};
test_label[4471] = '{32'h41357bc5};
test_output[4471] = '{32'h42a0ac0b};
/*############ DEBUG ############
test_input[35768:35775] = '{1.08577242916, 91.6787385721, 21.8712412228, 11.3427174274, 3.90077128115, -44.006394602, -3.56467593792, 16.3532903473};
test_label[4471] = '{11.3427174274};
test_output[4471] = '{80.3360211447};
############ END DEBUG ############*/
test_input[35776:35783] = '{32'h425291f0, 32'h40599433, 32'h411d27cc, 32'hc2018407, 32'h3fa1969f, 32'hc2ae4841, 32'h42b12515, 32'hc18f8890};
test_label[4472] = '{32'hc2ae4841};
test_output[4472] = '{32'h432fb6ab};
/*############ DEBUG ############
test_input[35776:35783] = '{52.6425160773, 3.39967035849, 9.8222157529, -32.3789331464, 1.26240907116, -87.1411171354, 88.5724256347, -17.9416814017};
test_label[4472] = '{-87.1411171354};
test_output[4472] = '{175.71354277};
############ END DEBUG ############*/
test_input[35784:35791] = '{32'h423118e2, 32'h429298a2, 32'h4273ef63, 32'h42b9b435, 32'hc19f4281, 32'h42a18055, 32'h428caa09, 32'hc2491d28};
test_label[4473] = '{32'hc2491d28};
test_output[4473] = '{32'h430f2165};
/*############ DEBUG ############
test_input[35784:35791] = '{44.2742992699, 73.2981147544, 60.983775739, 92.8519680411, -19.9074731756, 80.7506504834, 70.3321028638, -50.2784726519};
test_label[4473] = '{-50.2784726519};
test_output[4473] = '{143.130446249};
############ END DEBUG ############*/
test_input[35792:35799] = '{32'h41c07a60, 32'h42a3b049, 32'h42c69551, 32'h42b919d8, 32'hc2c46d43, 32'hc24d2ee2, 32'h4216a1f0, 32'h42349c60};
test_label[4474] = '{32'h42b919d8};
test_output[4474] = '{32'h40d7c145};
/*############ DEBUG ############
test_input[35792:35799] = '{24.0597527361, 81.8443051342, 99.2916361953, 92.5504741568, -98.2134030223, -51.2957828327, 37.6581402496, 45.152709834};
test_label[4474] = '{92.5504741568};
test_output[4474] = '{6.74234264146};
############ END DEBUG ############*/
test_input[35800:35807] = '{32'hc1be386f, 32'hc2b6e36f, 32'h405c226d, 32'h418a9a8e, 32'h42c66e4d, 32'h41bee431, 32'h42a253e1, 32'hc28fe582};
test_label[4475] = '{32'h42a253e1};
test_output[4475] = '{32'h419069b0};
/*############ DEBUG ############
test_input[35800:35807] = '{-23.7775554221, -91.4442080245, 3.43960111239, 17.325467033, 99.215434918, 23.8614211466, 81.1638295899, -71.9482610539};
test_label[4475] = '{81.1638295899};
test_output[4475] = '{18.0516053426};
############ END DEBUG ############*/
test_input[35808:35815] = '{32'h42a7ff94, 32'hc1e63499, 32'hc2c37b34, 32'hc2057402, 32'hc2b8966a, 32'h420ef0d1, 32'hc213c3e3, 32'hc229c0b0};
test_label[4476] = '{32'hc1e63499};
test_output[4476] = '{32'h42e18cbb};
/*############ DEBUG ############
test_input[35808:35815] = '{83.9991779591, -28.7756826754, -97.7406275308, -33.363289704, -92.2937795884, 35.7351733884, -36.9412966186, -42.4381726163};
test_label[4476] = '{-28.7756826754};
test_output[4476] = '{112.774860635};
############ END DEBUG ############*/
test_input[35816:35823] = '{32'hc08c7d08, 32'h428315b6, 32'h42a590c7, 32'hc180f03b, 32'hc216890a, 32'h428fd123, 32'hc269b0ce, 32'hc1c47686};
test_label[4477] = '{32'hc216890a};
test_output[4477] = '{32'h42f0d54f};
/*############ DEBUG ############
test_input[35816:35823] = '{-4.39026265339, 65.5424029798, 82.7827713704, -16.1172999075, -37.6338274878, 71.9084688241, -58.4226623569, -24.5578721195};
test_label[4477] = '{-37.6338274878};
test_output[4477] = '{120.416617829};
############ END DEBUG ############*/
test_input[35824:35831] = '{32'hc28603d5, 32'h426627c5, 32'h429c0325, 32'h42a0a6a7, 32'hc287a01a, 32'h4267fa07, 32'h4280d832, 32'h40871e1c};
test_label[4478] = '{32'h42a0a6a7};
test_output[4478] = '{32'h3dc01901};
/*############ DEBUG ############
test_input[35824:35831] = '{-67.007482889, 57.5388358847, 78.0061424045, 80.3254932818, -67.8127013281, 57.9941672741, 64.4222566259, 4.22242542153};
test_label[4478] = '{80.3254932818};
test_output[4478] = '{0.0937976931382};
############ END DEBUG ############*/
test_input[35832:35839] = '{32'h429f1926, 32'h42c0176c, 32'hc1cc5570, 32'h4229143f, 32'hc28c94c9, 32'hc184a500, 32'h41a12ab4, 32'hc225787d};
test_label[4479] = '{32'h42c0176c};
test_output[4479] = '{32'h339312c2};
/*############ DEBUG ############
test_input[35832:35839] = '{79.5491172381, 96.0457488492, -25.5417179724, 42.2697705111, -70.2905955388, -16.5805664633, 20.145852088, -41.3676629216};
test_label[4479] = '{96.0457488492};
test_output[4479] = '{6.84863319526e-08};
############ END DEBUG ############*/
test_input[35840:35847] = '{32'hc2498161, 32'hc2816e2d, 32'h428c9951, 32'hc1c470f2, 32'hc235408c, 32'hc189a9bd, 32'h42aed260, 32'hbfefb924};
test_label[4480] = '{32'hc235408c};
test_output[4480] = '{32'h4304b953};
/*############ DEBUG ############
test_input[35840:35847] = '{-50.3763457194, -64.7151855297, 70.2994449796, -24.5551490739, -45.3130322534, -17.2078804592, 87.410886323, -1.87283754788};
test_label[4480] = '{-45.3130322534};
test_output[4480] = '{132.723918613};
############ END DEBUG ############*/
test_input[35848:35855] = '{32'h4278b2c2, 32'hc1fa91af, 32'hc2afc745, 32'h42ba0a3d, 32'h42c4def3, 32'h428fb304, 32'h426d16fe, 32'h423d64ea};
test_label[4481] = '{32'hc1fa91af};
test_output[4481] = '{32'h4301c2d2};
/*############ DEBUG ############
test_input[35848:35855] = '{62.1745667326, -31.3211353582, -87.8892005509, 93.0200000913, 98.4354448268, 71.8496380467, 59.272454758, 47.3485488114};
test_label[4481] = '{-31.3211353582};
test_output[4481] = '{129.761017684};
############ END DEBUG ############*/
test_input[35856:35863] = '{32'hc242761f, 32'h42a225ee, 32'hc221d613, 32'h4180547d, 32'h41a78888, 32'h423cd1ae, 32'h41c2b488, 32'hc28993ad};
test_label[4482] = '{32'hc28993ad};
test_output[4482] = '{32'h4315dcce};
/*############ DEBUG ############
test_input[35856:35863] = '{-48.615351094, 81.0740851568, -40.4590549807, 16.0412538794, 20.9416661932, 47.204764159, 24.3381493576, -68.78843107};
test_label[4482] = '{-68.78843107};
test_output[4482] = '{149.862516227};
############ END DEBUG ############*/
test_input[35864:35871] = '{32'hc0ab94ff, 32'h428bb721, 32'hc266d7e5, 32'h42aa341e, 32'hc2179339, 32'h42a857f5, 32'hc2728476, 32'hc2c128ee};
test_label[4483] = '{32'h428bb721};
test_output[4483] = '{32'h41793a1e};
/*############ DEBUG ############
test_input[35864:35871] = '{-5.36193815084, 69.8576758022, -57.7108336018, 85.1017888563, -37.8937705043, 84.1717916825, -60.6293561355, -96.5799414228};
test_label[4483] = '{69.8576758022};
test_output[4483] = '{15.5766884687};
############ END DEBUG ############*/
test_input[35872:35879] = '{32'hc248c7a0, 32'h42a11db2, 32'h422deb2c, 32'h4093c351, 32'h41789b1a, 32'h42abac9f, 32'h4219ccdd, 32'h428c09fd};
test_label[4484] = '{32'h4219ccdd};
test_output[4484] = '{32'h423d9195};
/*############ DEBUG ############
test_input[35872:35879] = '{-50.1949465864, 80.5580010696, 43.4796613639, 4.61759238199, 15.5378669448, 85.8371478956, 38.4500617273, 70.0195049063};
test_label[4484] = '{38.4500617273};
test_output[4484] = '{47.3921701355};
############ END DEBUG ############*/
test_input[35880:35887] = '{32'h41e25425, 32'h42476c7c, 32'h426d9d58, 32'hc10a74f7, 32'h42ad2173, 32'hbe1636f3, 32'h425751f5, 32'hc21edee5};
test_label[4485] = '{32'h425751f5};
test_output[4485] = '{32'h4202f0f2};
/*############ DEBUG ############
test_input[35880:35887] = '{28.2910862325, 49.8559431239, 59.4036542942, -8.65355609899, 86.5653324839, -0.14669398449, 53.8300356411, -39.717669199};
test_label[4485] = '{53.8300356411};
test_output[4485] = '{32.7352968428};
############ END DEBUG ############*/
test_input[35888:35895] = '{32'h426a82bd, 32'hc2919efa, 32'h41f51f77, 32'h41e82138, 32'hc22bf24e, 32'h422bbd85, 32'hc25b1540, 32'h4187edcb};
test_label[4486] = '{32'h422bbd85};
test_output[4486] = '{32'h417b14e1};
/*############ DEBUG ############
test_input[35888:35895] = '{58.627673406, -72.8105038079, 30.6403628176, 29.016219787, -42.9866271227, 42.9350759072, -54.7707517578, 16.991110675};
test_label[4486] = '{42.9350759072};
test_output[4486] = '{15.6925976518};
############ END DEBUG ############*/
test_input[35896:35903] = '{32'hc2826057, 32'h421c99fb, 32'hc15e9d0a, 32'hc0393f4a, 32'hc261aa78, 32'h4139ca81, 32'h41f494ca, 32'h42143e98};
test_label[4487] = '{32'h421c99fb};
test_output[4487] = '{32'h3def5790};
/*############ DEBUG ############
test_input[35896:35903] = '{-65.1881609204, 39.1503703542, -13.9133392795, -2.89448796377, -56.4164738592, 11.6119397336, 30.5726508747, 37.0611274683};
test_label[4487] = '{39.1503703542};
test_output[4487] = '{0.116866233625};
############ END DEBUG ############*/
test_input[35904:35911] = '{32'h42bd79b5, 32'hc00a16e9, 32'h42b63b70, 32'h42690fe2, 32'hc2862467, 32'h4165b209, 32'h40a24734, 32'h422622a2};
test_label[4488] = '{32'h42bd79b5};
test_output[4488] = '{32'h3cd82c24};
/*############ DEBUG ############
test_input[35904:35911] = '{94.7377060922, -2.15764831668, 91.1160922003, 58.2655089029, -67.0710991037, 14.3559651571, 5.07119187606, 41.5338196665};
test_label[4488] = '{94.7377060922};
test_output[4488] = '{0.0263882347083};
############ END DEBUG ############*/
test_input[35912:35919] = '{32'h42300537, 32'hc264b32d, 32'h4115cd98, 32'hbce09c6e, 32'hc2b40fec, 32'h4286ee68, 32'hc2b0822e, 32'h4207e0dc};
test_label[4489] = '{32'h4115cd98};
test_output[4489] = '{32'h4268696a};
/*############ DEBUG ############
test_input[35912:35919] = '{44.0050929611, -57.1749765105, 9.36269376521, -0.0274183422804, -90.0310944339, 67.4656376107, -88.2542540135, 33.9695877116};
test_label[4489] = '{9.36269376521};
test_output[4489] = '{58.1029438455};
############ END DEBUG ############*/
test_input[35920:35927] = '{32'hc220ad56, 32'hc2447163, 32'hbf952ec0, 32'h4191c19d, 32'h425fee4d, 32'h42719b3d, 32'hc20bee27, 32'hc249250b};
test_label[4490] = '{32'h425fee4d};
test_output[4490] = '{32'h408dc996};
/*############ DEBUG ############
test_input[35920:35927] = '{-40.1692734405, -49.1107296401, -1.16548922173, 18.2195385199, 55.982717361, 60.401599478, -34.9825721524, -50.2861755689};
test_label[4490] = '{55.982717361};
test_output[4490] = '{4.43085781392};
############ END DEBUG ############*/
test_input[35928:35935] = '{32'hc239342f, 32'h42aab881, 32'hc266201d, 32'h421294d4, 32'h4295b296, 32'h4183a927, 32'hc27b6b62, 32'h40bf60a1};
test_label[4491] = '{32'h4295b296};
test_output[4491] = '{32'h41282f6e};
/*############ DEBUG ############
test_input[35928:35935] = '{-46.3009612985, 85.3603554469, -57.5313611761, 36.6453395238, 74.8488033429, 16.4575947771, -62.8548673334, 5.9805455903};
test_label[4491] = '{74.8488033429};
test_output[4491] = '{10.5115793239};
############ END DEBUG ############*/
test_input[35936:35943] = '{32'h42103f9e, 32'hc1b5ae3c, 32'h42a04d4c, 32'hc260f15c, 32'h4297bf8a, 32'hc2a7801b, 32'hc105a814, 32'hc20d8fb0};
test_label[4492] = '{32'h42103f9e};
test_output[4492] = '{32'h42306919};
/*############ DEBUG ############
test_input[35936:35943] = '{36.0621280111, -22.7100757826, 80.1509728786, -56.235702501, 75.8741022965, -83.75020926, -8.35353448157, -35.3903207291};
test_label[4492] = '{36.0621280111};
test_output[4492] = '{44.102635389};
############ END DEBUG ############*/
test_input[35944:35951] = '{32'h41a24441, 32'h424bc416, 32'h40a35bc8, 32'h428af58a, 32'h41476bcf, 32'hc20a7cc7, 32'h42b83066, 32'hc2b41f12};
test_label[4493] = '{32'h41476bcf};
test_output[4493] = '{32'h429f42ec};
/*############ DEBUG ############
test_input[35944:35951] = '{20.2833263238, 50.9414901178, 5.10495369162, 69.4795686899, 12.4638209254, -34.6218515316, 92.0945309488, -90.0606843246};
test_label[4493] = '{12.4638209254};
test_output[4493] = '{79.6307100236};
############ END DEBUG ############*/
test_input[35952:35959] = '{32'h42a043c0, 32'hc2c78de8, 32'hc18fa3e2, 32'h4242bad9, 32'hc29b1895, 32'hc217d58b, 32'hc1e24c5c, 32'h418c51d1};
test_label[4494] = '{32'hc217d58b};
test_output[4494] = '{32'h42ec2e85};
/*############ DEBUG ############
test_input[35952:35959] = '{80.1323231511, -99.7771596258, -17.9550215079, 48.6824675237, -77.5480100537, -37.9585390811, -28.2872852907, 17.5399495846};
test_label[4494] = '{-37.9585390811};
test_output[4494] = '{118.090862232};
############ END DEBUG ############*/
test_input[35960:35967] = '{32'hc250b77c, 32'h420bd035, 32'h428a51e0, 32'h40aff626, 32'hc2bfb77e, 32'hc2b16108, 32'hc249e167, 32'h428563a8};
test_label[4495] = '{32'h428563a8};
test_output[4495] = '{32'h4022ff61};
/*############ DEBUG ############
test_input[35960:35967] = '{-52.1791839096, 34.9533280171, 69.1599095891, 5.49879732684, -95.8583846912, -88.6895143298, -50.4701198822, 66.6946393549};
test_label[4495] = '{66.6946393549};
test_output[4495] = '{2.54683720097};
############ END DEBUG ############*/
test_input[35968:35975] = '{32'hc2b2fc65, 32'h41e9621c, 32'h4231c2f0, 32'h418a2228, 32'h42a81358, 32'h41a9ebd5, 32'hc203278d, 32'h423ea2d4};
test_label[4496] = '{32'h4231c2f0};
test_output[4496] = '{32'h421e63c0};
/*############ DEBUG ############
test_input[35968:35975] = '{-89.4929587833, 29.1729042696, 44.440369882, 17.2666777644, 84.0377814338, 21.2401526931, -32.7886257047, 47.6590102114};
test_label[4496] = '{44.440369882};
test_output[4496] = '{39.5974115518};
############ END DEBUG ############*/
test_input[35976:35983] = '{32'h41412216, 32'h42aec6d8, 32'hc29299ce, 32'hc2ad0156, 32'hc22b2530, 32'h428c60b1, 32'hc27e43fe, 32'h4295d39a};
test_label[4497] = '{32'h4295d39a};
test_output[4497] = '{32'h414799f9};
/*############ DEBUG ############
test_input[35976:35983] = '{12.0708218525, 87.3883699242, -73.3004025267, -86.5026080691, -42.7863161404, 70.1888506577, -63.5663985103, 74.9132828991};
test_label[4497] = '{74.9132828991};
test_output[4497] = '{12.4750908796};
############ END DEBUG ############*/
test_input[35984:35991] = '{32'hc03a648c, 32'hc2983c14, 32'h422f9eae, 32'hc18f8708, 32'hc231d928, 32'hc2676398, 32'hc1918e29, 32'h4179dd6f};
test_label[4498] = '{32'hc231d928};
test_output[4498] = '{32'h42b0bbeb};
/*############ DEBUG ############
test_input[35984:35991] = '{-2.91238696373, -76.1173408271, 43.90496129, -17.940933884, -44.4620648705, -57.8472583579, -18.1944133754, 15.6165607598};
test_label[4498] = '{-44.4620648705};
test_output[4498] = '{88.3670261605};
############ END DEBUG ############*/
test_input[35992:35999] = '{32'hc2a6d341, 32'hc223a694, 32'hc1e62867, 32'h42c7108e, 32'h4254dd8f, 32'hc2674433, 32'hc28ade7e, 32'h40b273ce};
test_label[4499] = '{32'h42c7108e};
test_output[4499] = '{32'h80000000};
/*############ DEBUG ############
test_input[35992:35999] = '{-83.4126078346, -40.9126751834, -28.7697272957, 99.5323330092, 53.2163644035, -57.8166010713, -69.4345533554, 5.57663627516};
test_label[4499] = '{99.5323330092};
test_output[4499] = '{-0.0};
############ END DEBUG ############*/
test_input[36000:36007] = '{32'h4265f41a, 32'h41024cc2, 32'h412dea65, 32'hc262eefb, 32'hc2379913, 32'hc223755f, 32'hc1f79ca7, 32'hc288f8c7};
test_label[4500] = '{32'hc223755f};
test_output[4500] = '{32'h42c4b4bc};
/*############ DEBUG ############
test_input[36000:36007] = '{57.488379317, 8.1437393169, 10.8697256965, -56.7333787206, -45.8994872872, -40.8646187773, -30.9514903183, -68.4858917711};
test_label[4500] = '{-40.8646187773};
test_output[4500] = '{98.3529980943};
############ END DEBUG ############*/
test_input[36008:36015] = '{32'hc1e45a5f, 32'hc24b94c2, 32'hc21aec0a, 32'h41d541ce, 32'h42807a08, 32'h4287ca33, 32'h427efb60, 32'hc282a3ee};
test_label[4501] = '{32'hc21aec0a};
test_output[4501] = '{32'h42d55515};
/*############ DEBUG ############
test_input[36008:36015] = '{-28.544125733, -50.8952729754, -38.7305079245, 26.6571303151, 64.2383436877, 67.8949182902, 63.7454832146, -65.320173309};
test_label[4501] = '{-38.7305079245};
test_output[4501] = '{106.666178574};
############ END DEBUG ############*/
test_input[36016:36023] = '{32'hc2860e87, 32'hc29e6d7b, 32'h42c1861b, 32'hc29e6eef, 32'h4231c3a8, 32'h42a8ea92, 32'hc21c41a0, 32'h4297e60c};
test_label[4502] = '{32'h42a8ea92};
test_output[4502] = '{32'h4144dc4a};
/*############ DEBUG ############
test_input[36016:36023] = '{-67.0283730702, -79.2138304889, 96.7619223155, -79.216667653, 44.4410689946, 84.458145139, -39.0640886325, 75.9493110636};
test_label[4502] = '{84.458145139};
test_output[4502] = '{12.3037817119};
############ END DEBUG ############*/
test_input[36024:36031] = '{32'h42843f90, 32'hc1965cb1, 32'h4239eb80, 32'hc2b9f447, 32'hc2602583, 32'hc234ee3a, 32'h4299c409, 32'hc244fcd5};
test_label[4503] = '{32'hc2b9f447};
test_output[4503] = '{32'h4329dc29};
/*############ DEBUG ############
test_input[36024:36031] = '{66.1241451169, -18.7952589342, 46.4799801094, -92.9771043636, -56.0366313894, -45.2326440177, 76.8828776099, -49.2469066147};
test_label[4503] = '{-92.9771043636};
test_output[4503] = '{169.860003232};
############ END DEBUG ############*/
test_input[36032:36039] = '{32'hc0b3479d, 32'h41ed8aab, 32'hbe92fe74, 32'h42696063, 32'h4280cde2, 32'h42165a36, 32'h405a44df, 32'h42c5750f};
test_label[4504] = '{32'hbe92fe74};
test_output[4504] = '{32'h42c6080e};
/*############ DEBUG ############
test_input[36032:36039] = '{-5.60249176731, 29.6927089781, -0.287097575461, 58.3441276334, 64.4021166093, 37.588096534, 3.41045350746, 98.72863268};
test_label[4504] = '{-0.287097575461};
test_output[4504] = '{99.0157302554};
############ END DEBUG ############*/
test_input[36040:36047] = '{32'hc2ba72d4, 32'hc262b3f6, 32'hc28c4d38, 32'h42193d27, 32'h429505df, 32'h41bda9d5, 32'hc2c52e33, 32'hc26f5ad2};
test_label[4505] = '{32'hc26f5ad2};
test_output[4505] = '{32'h430659a4};
/*############ DEBUG ############
test_input[36040:36047] = '{-93.2242714311, -56.6757440501, -70.1508211442, 38.3097172096, 74.5114637449, 23.7079251743, -98.5902315148, -59.8386927174};
test_label[4505] = '{-59.8386927174};
test_output[4505] = '{134.350156462};
############ END DEBUG ############*/
test_input[36048:36055] = '{32'hc1d608aa, 32'hc29ca4d7, 32'hc2bf5061, 32'h42a45014, 32'hc2349b58, 32'hc268cfd8, 32'h42c733f1, 32'h41806688};
test_label[4506] = '{32'hc2bf5061};
test_output[4506] = '{32'h43434229};
/*############ DEBUG ############
test_input[36048:36055] = '{-26.7542308033, -78.321949825, -95.6569880545, 82.1564055517, -45.1517035272, -58.2029742699, 99.6014487341, 16.0500645835};
test_label[4506] = '{-95.6569880545};
test_output[4506] = '{195.258436815};
############ END DEBUG ############*/
test_input[36056:36063] = '{32'h42b972ef, 32'hc249a2fc, 32'h4270a8de, 32'h42994da6, 32'h4129be7f, 32'hc275e6e3, 32'h42b28c77, 32'h42365950};
test_label[4507] = '{32'h42b972ef};
test_output[4507] = '{32'h3cfffc60};
/*############ DEBUG ############
test_input[36056:36063] = '{92.7244782683, -50.4091656828, 60.1649083036, 76.6516558259, 10.6090080279, -61.4754742623, 89.2743486056, 45.5872195753};
test_label[4507] = '{92.7244782683};
test_output[4507] = '{0.0312482723912};
############ END DEBUG ############*/
test_input[36064:36071] = '{32'hc2b6d864, 32'hc28612f5, 32'hc2885222, 32'hc230688d, 32'hc253c825, 32'hc1af5309, 32'hc29f2dfc, 32'h42b8804c};
test_label[4508] = '{32'hc29f2dfc};
test_output[4508] = '{32'h432bd724};
/*############ DEBUG ############
test_input[36064:36071] = '{-91.4226375283, -67.0370264034, -68.1604124366, -44.1020996762, -52.9454529943, -21.9155447188, -79.5898155207, 92.2505832486};
test_label[4508] = '{-79.5898155207};
test_output[4508] = '{171.840398769};
############ END DEBUG ############*/
test_input[36072:36079] = '{32'hc288967b, 32'hc2bc65ae, 32'h42a210cd, 32'h42227037, 32'h429dde09, 32'h41aeeede, 32'hc29211fb, 32'h41a66d25};
test_label[4509] = '{32'hc288967b};
test_output[4509] = '{32'h4315713c};
/*############ DEBUG ############
test_input[36072:36079] = '{-68.2939035608, -94.1985929759, 81.0328109574, 40.6095838422, 78.9336590397, 21.8666338316, -73.035119159, 20.8032930265};
test_label[4509] = '{-68.2939035608};
test_output[4509] = '{149.442326599};
############ END DEBUG ############*/
test_input[36080:36087] = '{32'hc2317000, 32'hc2b3c37f, 32'h42133f75, 32'hc202f020, 32'hc294c029, 32'hc29ded55, 32'h42c2cada, 32'hc236488c};
test_label[4510] = '{32'hc29ded55};
test_output[4510] = '{32'h43305c17};
/*############ DEBUG ############
test_input[36080:36087] = '{-44.3593757865, -89.881825429, 36.811971085, -32.7344982286, -74.3753143974, -78.963537126, 97.3961916274, -45.5708483561};
test_label[4510] = '{-78.963537126};
test_output[4510] = '{176.359728753};
############ END DEBUG ############*/
test_input[36088:36095] = '{32'hc2085371, 32'h429ab6d9, 32'h424a2a26, 32'h4064bbdd, 32'hc29be780, 32'hc19b132a, 32'hc1ff49e2, 32'h42a9287d};
test_label[4511] = '{32'h424a2a26};
test_output[4511] = '{32'h42082793};
/*############ DEBUG ############
test_input[36088:36095] = '{-34.08148559, 77.3571273998, 50.5411612969, 3.57396619911, -77.9521461973, -19.3843569164, -31.9110752227, 84.5790769003};
test_label[4511] = '{50.5411612969};
test_output[4511] = '{34.038645714};
############ END DEBUG ############*/
test_input[36096:36103] = '{32'hc2bf6232, 32'h42835cc5, 32'hc26554f4, 32'h4299d15c, 32'h423fb516, 32'hc297497d, 32'hc1621fe6, 32'hc26d29b5};
test_label[4512] = '{32'h42835cc5};
test_output[4512] = '{32'h4133a4c9};
/*############ DEBUG ############
test_input[36096:36103] = '{-95.6917898968, 65.6811892176, -57.3329613529, 76.9089063478, 47.9268421122, -75.6435295816, -14.1327872831, -59.2907295104};
test_label[4512] = '{65.6811892176};
test_output[4512] = '{11.2277304305};
############ END DEBUG ############*/
test_input[36104:36111] = '{32'h426aa601, 32'h424fd9f6, 32'hc22427b2, 32'hc21f496b, 32'h422da63d, 32'hc2bf8d37, 32'h428b5d3b, 32'h40c81ea2};
test_label[4513] = '{32'h426aa601};
test_output[4513] = '{32'h413051e6};
/*############ DEBUG ############
test_input[36104:36111] = '{58.6621115453, 51.9628519309, -41.0387663164, -39.8216983617, 43.4123428031, -95.7758109256, 69.6820898449, 6.2537395021};
test_label[4513] = '{58.6621115453};
test_output[4513] = '{11.019994691};
############ END DEBUG ############*/
test_input[36112:36119] = '{32'h41de9d2d, 32'hc0289a6e, 32'hc29369b6, 32'hc20d46ac, 32'hc28a5145, 32'hc278188c, 32'hc1af4a21, 32'h4223a683};
test_label[4514] = '{32'hc0289a6e};
test_output[4514] = '{32'h422e302b};
/*############ DEBUG ############
test_input[36112:36119] = '{27.8267452974, -2.63442563314, -73.7064656522, -35.3190144834, -69.1587260697, -62.0239703411, -21.9111949987, 40.9126103797};
test_label[4514] = '{-2.63442563314};
test_output[4514] = '{43.5470380872};
############ END DEBUG ############*/
test_input[36120:36127] = '{32'h429bc20e, 32'h42c66dd5, 32'hc1937a1a, 32'hc2c626ba, 32'hc2bcc94a, 32'hc180befc, 32'h42b12956, 32'hc29951b9};
test_label[4515] = '{32'hc2bcc94a};
test_output[4515] = '{32'h43419b91};
/*############ DEBUG ############
test_input[36120:36127] = '{77.8790102618, 99.2145154003, -18.4346192933, -99.0756389967, -94.3931399085, -16.0932531633, 88.5807319677, -76.6596138324};
test_label[4515] = '{-94.3931399085};
test_output[4515] = '{193.607679397};
############ END DEBUG ############*/
test_input[36128:36135] = '{32'h4206b7e7, 32'hc29f1d86, 32'h41e6b383, 32'h40870f3b, 32'hc21e35b9, 32'h423fe9b2, 32'h42b0136b, 32'h427e0ffd};
test_label[4516] = '{32'h4206b7e7};
test_output[4516] = '{32'h42596ef0};
/*############ DEBUG ############
test_input[36128:36135] = '{33.6795928022, -79.5576601406, 28.83765195, 4.22060904773, -39.5524643787, 47.9782193049, 88.0379286734, 63.5156140697};
test_label[4516] = '{33.6795928022};
test_output[4516] = '{54.3583358713};
############ END DEBUG ############*/
test_input[36136:36143] = '{32'hc2b08a7d, 32'h4296274c, 32'h41dc9a0e, 32'h420b137e, 32'hc03daa34, 32'hc23de5d0, 32'h40728ca3, 32'hc27d727d};
test_label[4517] = '{32'h4296274c};
test_output[4517] = '{32'h80000000};
/*############ DEBUG ############
test_input[36136:36143] = '{-88.2704849467, 75.0767549464, 27.5752218806, 34.7690344557, -2.96351328093, -47.4744274887, 3.78983375243, -63.3618061777};
test_label[4517] = '{75.0767549464};
test_output[4517] = '{-0.0};
############ END DEBUG ############*/
test_input[36144:36151] = '{32'hc2882943, 32'hc2290bfe, 32'hc2481e35, 32'hc21d0160, 32'hc145588b, 32'h4186c87d, 32'h4213cc01, 32'hc2304387};
test_label[4518] = '{32'hc2290bfe};
test_output[4518] = '{32'h429e6bff};
/*############ DEBUG ############
test_input[36144:36151] = '{-68.0805860334, -42.2617111995, -50.0294974471, -39.251341048, -12.3341170833, 16.8478954543, 36.9492208446, -44.0659445275};
test_label[4518] = '{-42.2617111995};
test_output[4518] = '{79.210932046};
############ END DEBUG ############*/
test_input[36152:36159] = '{32'hc0a05ab7, 32'h4197a297, 32'hc1bbbee8, 32'h41f3d4e0, 32'hbfd1e355, 32'hc1f6578a, 32'h422a9135, 32'hc1713dbe};
test_label[4519] = '{32'hbfd1e355};
test_output[4519] = '{32'h42312051};
/*############ DEBUG ############
test_input[36152:36159] = '{-5.01107376746, 18.954389057, -23.4682167687, 30.4789424283, -1.63975013733, -30.7927436391, 42.641803303, -15.0775735885};
test_label[4519] = '{-1.63975013733};
test_output[4519] = '{44.2815586612};
############ END DEBUG ############*/
test_input[36160:36167] = '{32'hc2ba4476, 32'hc2ab031a, 32'hc2b2a6f0, 32'h42839026, 32'hc2aadf3a, 32'h42b8b417, 32'hc290e28d, 32'hc1470f9e};
test_label[4520] = '{32'hc1470f9e};
test_output[4520] = '{32'h42d1960b};
/*############ DEBUG ############
test_input[36160:36167] = '{-93.1337136904, -85.5060558733, -89.3260491537, 65.7815432299, -85.4359929465, 92.3517382066, -72.4424810858, -12.4413132609};
test_label[4520] = '{-12.4413132609};
test_output[4520] = '{104.793051467};
############ END DEBUG ############*/
test_input[36168:36175] = '{32'h4282d53f, 32'hc263a272, 32'hc16a966a, 32'h428efb24, 32'h428c8a32, 32'hc1118ed3, 32'hc225e9e8, 32'h42c0d43e};
test_label[4521] = '{32'hc1118ed3};
test_output[4521] = '{32'h42d30618};
/*############ DEBUG ############
test_input[36168:36175] = '{65.4164977934, -56.9086386756, -14.6617224752, 71.4905120834, 70.2699135559, -9.09736877738, -41.4784222289, 96.414536737};
test_label[4521] = '{-9.09736877738};
test_output[4521] = '{105.511905514};
############ END DEBUG ############*/
test_input[36176:36183] = '{32'hc2a34827, 32'h42ad5c27, 32'h410c7638, 32'hc1c8f781, 32'hc284226b, 32'hc1ea62cb, 32'hc286a85c, 32'h42374aef};
test_label[4522] = '{32'hc286a85c};
test_output[4522] = '{32'h431a0242};
/*############ DEBUG ############
test_input[36176:36183] = '{-81.6409199571, 86.6799868021, 8.77886232609, -25.1208522538, -66.0672214983, -29.2982382872, -67.328830604, 45.8231765061};
test_label[4522] = '{-67.328830604};
test_output[4522] = '{154.008817406};
############ END DEBUG ############*/
test_input[36184:36191] = '{32'h429d70d1, 32'hc2450d6b, 32'hc2105df4, 32'h42bc36c6, 32'hc1e35005, 32'h42c7d2c2, 32'hc25c95a4, 32'hc26f2794};
test_label[4523] = '{32'h42bc36c6};
test_output[4523] = '{32'h40b9d872};
/*############ DEBUG ############
test_input[36184:36191] = '{78.7203431637, -49.2631027633, -36.0917522328, 94.1069763352, -28.4140712589, 99.9116390449, -55.146132278, -59.7886497524};
test_label[4523] = '{94.1069763352};
test_output[4523] = '{5.80767164998};
############ END DEBUG ############*/
test_input[36192:36199] = '{32'hc2aa3f41, 32'h42285877, 32'hc2725d65, 32'hc220f89c, 32'hc11cfcb8, 32'h42967180, 32'hc2b9dd0f, 32'h420fe83b};
test_label[4524] = '{32'h42967180};
test_output[4524] = '{32'h27900000};
/*############ DEBUG ############
test_input[36192:36199] = '{-85.1235400956, 42.0863919527, -60.5912059326, -40.2427820799, -9.81169901186, 75.2216822878, -92.9317541478, 35.9767892293};
test_label[4524] = '{75.2216822878};
test_output[4524] = '{3.99680288865e-15};
############ END DEBUG ############*/
test_input[36200:36207] = '{32'h4249fb0c, 32'h420d2947, 32'hc0ece446, 32'hc27e1334, 32'hc2892027, 32'hc0b711d9, 32'h418e2d1f, 32'hc25ba263};
test_label[4525] = '{32'h4249fb0c};
test_output[4525] = '{32'h3485cf28};
/*############ DEBUG ############
test_input[36200:36207] = '{50.4951621062, 35.2903089579, -7.40286528195, -63.5187537473, -68.5628001803, -5.72092853004, 17.7720309663, -54.908582404};
test_label[4525] = '{50.4951621062};
test_output[4525] = '{2.49239078128e-07};
############ END DEBUG ############*/
test_input[36208:36215] = '{32'hc2b9e2de, 32'h42c212fc, 32'h42be0c66, 32'hc22e61a8, 32'h42032063, 32'hc10d2758, 32'h41a0bf9d, 32'hc19ef16e};
test_label[4526] = '{32'h42be0c66};
test_output[4526] = '{32'h4008d95c};
/*############ DEBUG ############
test_input[36208:36215] = '{-92.9430969208, 97.0370761111, 95.0242128789, -43.5953661323, 32.7816262307, -8.8221057259, 20.0935617138, -19.867885386};
test_label[4526] = '{95.0242128789};
test_output[4526] = '{2.13826656628};
############ END DEBUG ############*/
test_input[36216:36223] = '{32'hc1cb5b0d, 32'hc2b00fad, 32'hc2072a24, 32'hc204c4e1, 32'hc2a35d87, 32'h41d71c3c, 32'hc17ea192, 32'h41d6b501};
test_label[4527] = '{32'hc2072a24};
test_output[4527] = '{32'h4275648f};
/*############ DEBUG ############
test_input[36216:36223] = '{-25.4194575463, -88.0306159718, -33.7911523531, -33.192266454, -81.6826735492, 26.8887870752, -15.9144457903, 26.8383806504};
test_label[4527] = '{-33.7911523531};
test_output[4527] = '{61.3482009638};
############ END DEBUG ############*/
test_input[36224:36231] = '{32'hc237dc2c, 32'hc2676f38, 32'hc286b4f8, 32'h42b6361c, 32'hc2a979a3, 32'hc08d5197, 32'hc2a628bb, 32'h429375d5};
test_label[4528] = '{32'hc2a628bb};
test_output[4528] = '{32'h432e2f6c};
/*############ DEBUG ############
test_input[36224:36231] = '{-45.9650121849, -57.8586120696, -67.3534543781, 91.1056854198, -84.7375722952, -4.41620985275, -83.0795551441, 73.7301414408};
test_label[4528] = '{-83.0795551441};
test_output[4528] = '{174.185240592};
############ END DEBUG ############*/
test_input[36232:36239] = '{32'h41b38e62, 32'h42c5613d, 32'hc2a8e10c, 32'hc2229964, 32'h41e0b619, 32'hc2a16861, 32'h428ef9cb, 32'hc11482db};
test_label[4529] = '{32'hc2a8e10c};
test_output[4529] = '{32'h43372124};
/*############ DEBUG ############
test_input[36232:36239] = '{22.4445233426, 98.6899193899, -84.4395431371, -40.6497945725, 28.0889143763, -80.7038686697, 71.4878744297, -9.28194675737};
test_label[4529] = '{-84.4395431371};
test_output[4529] = '{183.129462527};
############ END DEBUG ############*/
test_input[36240:36247] = '{32'h42a8f8ea, 32'hc297b836, 32'h426ab2a7, 32'hc1a9f5b4, 32'hc1a4b978, 32'h4194bd32, 32'hc2934a02, 32'hc1c28f60};
test_label[4530] = '{32'hc2934a02};
test_output[4530] = '{32'h431e2176};
/*############ DEBUG ############
test_input[36240:36247] = '{84.4861609938, -75.8597833603, 58.6744637695, -21.2449727521, -20.5905607634, 18.5923807951, -73.6445445338, -24.3200081667};
test_label[4530] = '{-73.6445445338};
test_output[4530] = '{158.130705528};
############ END DEBUG ############*/
test_input[36248:36255] = '{32'h42299d27, 32'h419d5e8f, 32'h4273fd29, 32'hc0f778e6, 32'hbe25af12, 32'h41baa95f, 32'h42a9833b, 32'h42528d53};
test_label[4531] = '{32'h41baa95f};
test_output[4531] = '{32'h4275b1c6};
/*############ DEBUG ############
test_input[36248:36255] = '{42.4034686684, 19.6711719525, 60.9972252725, -7.73350833496, -0.161800648762, 23.3327006117, 84.7563078784, 52.6380101258};
test_label[4531] = '{23.3327006117};
test_output[4531] = '{61.4236072668};
############ END DEBUG ############*/
test_input[36256:36263] = '{32'h4143878f, 32'h42949f2d, 32'hc20778f2, 32'hbed917af, 32'h41e7cea5, 32'h429f29af, 32'hc21e1295, 32'h42c4ee13};
test_label[4532] = '{32'h42949f2d};
test_output[4532] = '{32'h41c13b96};
/*############ DEBUG ############
test_input[36256:36263] = '{12.2205951018, 74.3108908175, -33.8681089678, -0.424008821408, 28.9759003332, 79.5814132197, -39.518148318, 98.4649862358};
test_label[4532] = '{74.3108908175};
test_output[4532] = '{24.1540954246};
############ END DEBUG ############*/
test_input[36264:36271] = '{32'hc1d7115f, 32'h42839984, 32'hc25c27c5, 32'hc2ab8984, 32'hc0215a65, 32'h4107c79f, 32'h41518b99, 32'hc27ed460};
test_label[4533] = '{32'hc0215a65};
test_output[4533] = '{32'h4288a457};
/*############ DEBUG ############
test_input[36264:36271] = '{-26.8834823546, 65.7998370939, -55.0388392818, -85.7685872615, -2.52114223862, 8.48623530329, 13.0965815069, -63.7073973655};
test_label[4533] = '{-2.52114223862};
test_output[4533] = '{68.3209793325};
############ END DEBUG ############*/
test_input[36272:36279] = '{32'hc0ed1d5c, 32'h42149d16, 32'hc1565047, 32'h42b27e8f, 32'h42687b82, 32'hc2562b02, 32'hc2b077e2, 32'h428a0c1a};
test_label[4534] = '{32'hc0ed1d5c};
test_output[4534] = '{32'h42c15065};
/*############ DEBUG ############
test_input[36272:36279] = '{-7.40983411654, 37.1534027852, -13.394598623, 89.2471877731, 58.1206113787, -53.5420008704, -88.2341496777, 69.023633173};
test_label[4534] = '{-7.40983411654};
test_output[4534] = '{96.6570218913};
############ END DEBUG ############*/
test_input[36280:36287] = '{32'h42397c94, 32'hc176262e, 32'h3ecb3a16, 32'hc29fbc94, 32'hc2ac0a0c, 32'hc25e52b2, 32'hc2abc7cb, 32'h41f0f673};
test_label[4535] = '{32'hc29fbc94};
test_output[4535] = '{32'h42fc7ade};
/*############ DEBUG ############
test_input[36280:36287] = '{46.3716574801, -15.384321289, 0.396927548706, -79.8683184183, -86.0196204068, -55.5807577162, -85.8902244165, 30.1203357235};
test_label[4535] = '{-79.8683184183};
test_output[4535] = '{126.239975986};
############ END DEBUG ############*/
test_input[36288:36295] = '{32'hc27277c4, 32'h42b7083d, 32'hc1f9c94c, 32'h426acdde, 32'h41a44b1d, 32'hc2c3ac78, 32'h422d0cb1, 32'hc1317e93};
test_label[4536] = '{32'h426acdde};
test_output[4536] = '{32'h4203429d};
/*############ DEBUG ############
test_input[36288:36295] = '{-60.616957427, 91.5160938744, -31.2232890386, 58.7010423491, 20.5366757392, -97.8368505752, 43.2623937353, -11.0934015452};
test_label[4536] = '{58.7010423491};
test_output[4536] = '{32.8150515253};
############ END DEBUG ############*/
test_input[36296:36303] = '{32'hc180a449, 32'hc1911ab5, 32'hc2857dd9, 32'h428f5084, 32'h42a35e06, 32'h42a2f55b, 32'hc20ce532, 32'h41c6f3bf};
test_label[4537] = '{32'hc2857dd9};
test_output[4537] = '{32'h4315068e};
/*############ DEBUG ############
test_input[36296:36303] = '{-16.0802164937, -18.1380413091, -66.7457980974, 71.6572600256, 81.6836415204, 81.4792075078, -35.2238222474, 24.8690167867};
test_label[4537] = '{-66.7457980974};
test_output[4537] = '{149.025609239};
############ END DEBUG ############*/
test_input[36304:36311] = '{32'h42419d10, 32'h4212a3c2, 32'h42bab7f3, 32'h42c57069, 32'hc0aebf87, 32'hc240a656, 32'hc209142c, 32'h42926f80};
test_label[4538] = '{32'h4212a3c2};
test_output[4538] = '{32'h427841dc};
/*############ DEBUG ############
test_input[36304:36311] = '{48.4033795236, 36.659919957, 93.3592769359, 98.7195485314, -5.46087960144, -48.1624365917, -34.2696995459, 73.2177708552};
test_label[4538] = '{36.659919957};
test_output[4538] = '{62.0643171952};
############ END DEBUG ############*/
test_input[36312:36319] = '{32'hc19c3db9, 32'hc27d30ce, 32'hc1e86940, 32'h41b59553, 32'h426f4bbe, 32'hc136339c, 32'hc24c259e, 32'h4267666a};
test_label[4539] = '{32'hc136339c};
test_output[4539] = '{32'h428eaeeb};
/*############ DEBUG ############
test_input[36312:36319] = '{-19.530138275, -63.2976625542, -29.0513911787, 22.6979113942, 59.8239660527, -11.3875997816, -51.036737026, 57.8500140007};
test_label[4539] = '{-11.3875997816};
test_output[4539] = '{71.341634692};
############ END DEBUG ############*/
test_input[36320:36327] = '{32'hc26cbb5e, 32'hc25c5802, 32'hc2ab0e20, 32'hc28eef81, 32'h42a6d90e, 32'h4269b057, 32'hc29afdec, 32'h42b92e47};
test_label[4540] = '{32'hc26cbb5e};
test_output[4540] = '{32'h4317c602};
/*############ DEBUG ############
test_input[36320:36327] = '{-59.1829740925, -55.0859440275, -85.5275890369, -71.4677814864, 83.423936796, 58.4222070693, -77.495941093, 92.5903860545};
test_label[4540] = '{-59.1829740925};
test_output[4540] = '{151.773464628};
############ END DEBUG ############*/
test_input[36328:36335] = '{32'h40ab5940, 32'h4292ac20, 32'hc1dcd5bc, 32'h42b48648, 32'h40b61470, 32'h41dcffff, 32'hc2961147, 32'h4262ab54};
test_label[4541] = '{32'h40ab5940};
test_output[4541] = '{32'h42a9d0b4};
/*############ DEBUG ############
test_input[36328:36335] = '{5.35464488056, 73.336181057, -27.6043628763, 90.2622698588, 5.68999471117, 27.6249980126, -75.0337434024, 56.6673136699};
test_label[4541] = '{5.35464488056};
test_output[4541] = '{84.9076250228};
############ END DEBUG ############*/
test_input[36336:36343] = '{32'hc273f261, 32'hc1fcbd56, 32'h429a35d6, 32'h429ad5ae, 32'h40ba7669, 32'hc1954c4f, 32'hc15e30f0, 32'hc233de07};
test_label[4542] = '{32'hc233de07};
test_output[4542] = '{32'h42f5dde1};
/*############ DEBUG ############
test_input[36336:36343] = '{-60.9866987625, -31.5924497399, 77.1051509928, 77.4173454135, 5.82695430665, -18.6622600545, -13.8869479216, -44.9668254074};
test_label[4542] = '{-44.9668254074};
test_output[4542] = '{122.933354803};
############ END DEBUG ############*/
test_input[36344:36351] = '{32'h4197ddd2, 32'hc29d038c, 32'hc29b20fd, 32'hc10740df, 32'h41179c7e, 32'h428d3e78, 32'h423c9f5c, 32'hc285bfa0};
test_label[4543] = '{32'hc29b20fd};
test_output[4543] = '{32'h43142fba};
/*############ DEBUG ############
test_input[36344:36351] = '{18.9833103588, -78.5069238728, -77.5644266766, -8.45333721212, 9.47570596089, 70.6220121768, 47.155625918, -66.8742711733};
test_label[4543] = '{-77.5644266766};
test_output[4543] = '{148.186438853};
############ END DEBUG ############*/
test_input[36352:36359] = '{32'h427741a8, 32'hc279627e, 32'hc1887844, 32'hc08f3dd0, 32'hc2127802, 32'h422f094d, 32'h42aad7e6, 32'hc146c612};
test_label[4544] = '{32'hc1887844};
test_output[4544] = '{32'h42ccf5f7};
/*############ DEBUG ############
test_input[36352:36359] = '{61.8141159814, -62.3461822321, -17.0587231167, -4.47629543733, -36.6171947168, 43.7590810403, 85.4216778023, -12.4233567949};
test_label[4544] = '{-17.0587231167};
test_output[4544] = '{102.480400919};
############ END DEBUG ############*/
test_input[36360:36367] = '{32'hc252abed, 32'h41f3dd2a, 32'hc1358bfc, 32'hc1acf509, 32'hc2034d50, 32'h42c5a4c2, 32'h40d6c837, 32'h42a8aae9};
test_label[4545] = '{32'h42c5a4c2};
test_output[4545] = '{32'h35090586};
/*############ DEBUG ############
test_input[36360:36367] = '{-52.6678976396, 30.4829909512, -11.3466763269, -21.6196467805, -32.8255015952, 98.82179409, 6.71194013074, 84.3338116558};
test_label[4545] = '{98.82179409};
test_output[4545] = '{5.10445129213e-07};
############ END DEBUG ############*/
test_input[36368:36375] = '{32'hc2c3e59f, 32'hc25ac8f5, 32'h420b3c0c, 32'hc2bb6e8d, 32'h423d5a98, 32'h4084dcd3, 32'h42477993, 32'hc29c00d8};
test_label[4546] = '{32'h42477993};
test_output[4546] = '{32'h3d9cee77};
/*############ DEBUG ############
test_input[36368:36375] = '{-97.9484821564, -54.6962470513, 34.80864017, -93.7159183046, 47.3384713729, 4.15195594975, 49.8687265836, -78.0016463797};
test_label[4546] = '{49.8687265836};
test_output[4546] = '{0.0766267085004};
############ END DEBUG ############*/
test_input[36376:36383] = '{32'hc20f889b, 32'h42120cb0, 32'hc27ddcdb, 32'h41a5a66c, 32'h4221ec57, 32'hc290e2e6, 32'hc28ff4c8, 32'h427d5fcd};
test_label[4547] = '{32'h42120cb0};
test_output[4547] = '{32'h41d6a63a};
/*############ DEBUG ############
test_input[36376:36383] = '{-35.8834024836, 36.5123904532, -63.4656792615, 20.7062608354, 40.4808007115, -72.4431616456, -71.9780920048, 63.3435566831};
test_label[4547] = '{36.5123904532};
test_output[4547] = '{26.83116623};
############ END DEBUG ############*/
test_input[36384:36391] = '{32'hc29051fb, 32'hc1b24702, 32'hc195c66d, 32'hc2a96541, 32'hc2ab05db, 32'hc0b493ed, 32'hc2616796, 32'hc29a323b};
test_label[4548] = '{32'hc2ab05db};
test_output[4548] = '{32'h429fbc9c};
/*############ DEBUG ############
test_input[36384:36391] = '{-72.160116097, -22.2846711349, -18.7218877412, -84.697762824, -85.5114355047, -5.64305732048, -56.3511566854, -77.0981090225};
test_label[4548] = '{-85.5114355047};
test_output[4548] = '{79.8683803325};
############ END DEBUG ############*/
test_input[36392:36399] = '{32'hc2b41f95, 32'hc29eda8e, 32'hc2bbcfdc, 32'h41a78fd7, 32'h42809992, 32'h4222e797, 32'hc29310f6, 32'hc2a46b1f};
test_label[4549] = '{32'h41a78fd7};
test_output[4549] = '{32'h422d6b38};
/*############ DEBUG ############
test_input[36392:36399] = '{-90.0616825959, -79.4268682209, -93.9059779895, 20.9452352391, 64.2999424744, 40.7261605179, -73.5331268755, -82.2092203796};
test_label[4549] = '{20.9452352391};
test_output[4549] = '{43.3547072354};
############ END DEBUG ############*/
test_input[36400:36407] = '{32'h42c1da62, 32'h428638fe, 32'hc29816ff, 32'hc2b93c67, 32'h41f0914b, 32'hc1f7b493, 32'hc1146f0e, 32'h414a1dfb};
test_label[4550] = '{32'hc29816ff};
test_output[4550] = '{32'h432cf8b0};
/*############ DEBUG ############
test_input[36400:36407] = '{96.9265286666, 67.1113158532, -76.0449122579, -92.617976703, 30.0709442427, -30.9631714625, -9.27711328829, 12.6323199024};
test_label[4550] = '{-76.0449122579};
test_output[4550] = '{172.971440925};
############ END DEBUG ############*/
test_input[36408:36415] = '{32'h41e1afa0, 32'hc24c0161, 32'h4208acf7, 32'hc24d6934, 32'h417f9bdd, 32'h42841c3e, 32'hc1ff2b15, 32'h42aeb889};
test_label[4551] = '{32'h4208acf7};
test_output[4551] = '{32'h4254c41b};
/*############ DEBUG ############
test_input[36408:36415] = '{28.2107547823, -51.00134749, 34.1689095124, -51.3527387478, 15.9755530275, 66.0551569086, -31.8960362873, 87.3604181592};
test_label[4551] = '{34.1689095124};
test_output[4551] = '{53.1915086473};
############ END DEBUG ############*/
test_input[36416:36423] = '{32'hc295e691, 32'h42117e78, 32'h425d974a, 32'hc221178d, 32'h41dbc48f, 32'hc2b4a025, 32'h413f3180, 32'hc23b5c06};
test_label[4552] = '{32'hc295e691};
test_output[4552] = '{32'h4302591b};
/*############ DEBUG ############
test_input[36416:36423] = '{-74.9503239474, 36.373505752, 55.3977420393, -40.2729977553, 27.4709760146, -90.3127790243, 11.9495847766, -46.8398651095};
test_label[4552] = '{-74.9503239474};
test_output[4552] = '{130.348065992};
############ END DEBUG ############*/
test_input[36424:36431] = '{32'hc1cb3471, 32'hc27d5ad1, 32'h424cbe47, 32'h423a1f4b, 32'hc2088a2d, 32'h42b938e3, 32'hc1cdf1bb, 32'hc1e151c1};
test_label[4553] = '{32'hc1cdf1bb};
test_output[4553] = '{32'h42ecb552};
/*############ DEBUG ############
test_input[36424:36431] = '{-25.4006060474, -63.3386875167, 51.185817796, 46.5305612427, -34.1349390176, 92.6111050675, -25.7430328896, -28.1649196138};
test_label[4553] = '{-25.7430328896};
test_output[4553] = '{118.354137957};
############ END DEBUG ############*/
test_input[36432:36439] = '{32'h425436d5, 32'h423814e0, 32'hc21a7eda, 32'hc28e9250, 32'hc28b2885, 32'hc27628f2, 32'hc29c22c2, 32'hc1e98769};
test_label[4554] = '{32'hc21a7eda};
test_output[4554] = '{32'h42b75b4b};
/*############ DEBUG ############
test_input[36432:36439] = '{53.0535467065, 46.0203855491, -38.6238795934, -71.2857653863, -69.5791433098, -61.5399858591, -78.0678863677, -29.1911187009};
test_label[4554] = '{-38.6238795934};
test_output[4554] = '{91.6783080498};
############ END DEBUG ############*/
test_input[36440:36447] = '{32'hc295b7c9, 32'hc206d9c7, 32'h418d0733, 32'hc2120be8, 32'h4234a7af, 32'h42c306fd, 32'h427b1e0b, 32'hc238a5fa};
test_label[4555] = '{32'hc206d9c7};
test_output[4555] = '{32'h430339f0};
/*############ DEBUG ############
test_input[36440:36447] = '{-74.8589574964, -33.7126738948, 17.6285159879, -36.5116259221, 45.1637541795, 97.5136472724, 62.7793391677, -46.1620853089};
test_label[4555] = '{-33.7126738948};
test_output[4555] = '{131.226321167};
############ END DEBUG ############*/
test_input[36448:36455] = '{32'h416a0721, 32'h41452a2a, 32'h429af02d, 32'h41978a01, 32'h3f2860f2, 32'hc2b4931c, 32'h424727ef, 32'h41609f96};
test_label[4556] = '{32'h416a0721};
test_output[4556] = '{32'h427b5e92};
/*############ DEBUG ############
test_input[36448:36455] = '{14.6267399873, 12.3227939954, 77.4690941096, 18.9423853301, 0.657729244031, -90.2873204145, 49.7889968228, 14.0389610329};
test_label[4556] = '{14.6267399873};
test_output[4556] = '{62.8423541223};
############ END DEBUG ############*/
test_input[36456:36463] = '{32'h422168e0, 32'hbfca08c5, 32'h42b7f496, 32'h42123d37, 32'h42906fc5, 32'h423e6744, 32'hc2671218, 32'hc27c5c5e};
test_label[4557] = '{32'h423e6744};
test_output[4557] = '{32'h423181e8};
/*############ DEBUG ############
test_input[36456:36463] = '{40.3524164206, -1.5783925677, 91.9777069874, 36.559778334, 72.2183013642, 47.6008460737, -57.7676709341, -63.0902018091};
test_label[4557] = '{47.6008460737};
test_output[4557] = '{44.3768609163};
############ END DEBUG ############*/
test_input[36464:36471] = '{32'hc2230211, 32'h41eb82f6, 32'hc29448c6, 32'hc2b61a46, 32'h42ace260, 32'hc259a9c5, 32'hc1cacfa2, 32'h42b4c495};
test_label[4558] = '{32'h42ace260};
test_output[4558] = '{32'h407d81aa};
/*############ DEBUG ############
test_input[36464:36471] = '{-40.7520195916, 29.4389465881, -74.1421321203, -91.0513178888, 86.4421375214, -54.4157914776, -25.3513826114, 90.3839496152};
test_label[4558] = '{86.4421375214};
test_output[4558] = '{3.96103906979};
############ END DEBUG ############*/
test_input[36472:36479] = '{32'h4076f28e, 32'h42a1796a, 32'h41f72b39, 32'h4267b00e, 32'h40c02076, 32'hc15008c7, 32'hbdab77d8, 32'h42aab428};
test_label[4559] = '{32'hbdab77d8};
test_output[4559] = '{32'h42aae412};
/*############ DEBUG ############
test_input[36472:36479] = '{3.85855435188, 80.7371362103, 30.8961054131, 57.9219276738, 6.00396273822, -13.0021428061, -0.0837246797182, 85.3518661155};
test_label[4559] = '{-0.0837246797182};
test_output[4559] = '{85.4454469219};
############ END DEBUG ############*/
test_input[36480:36487] = '{32'hc2ad327e, 32'hc29d5669, 32'hc2a0fd38, 32'hc2bfb658, 32'hc2706674, 32'h4294bfd7, 32'hc21b978d, 32'h429654d4};
test_label[4560] = '{32'hc2706674};
test_output[4560] = '{32'h4307a3bf};
/*############ DEBUG ############
test_input[36480:36487] = '{-86.5986213294, -78.6687682461, -80.4945669594, -95.856142735, -60.100053325, 74.3746899171, -38.8980003223, 75.1656829321};
test_label[4560] = '{-60.100053325};
test_output[4560] = '{135.639638005};
############ END DEBUG ############*/
test_input[36488:36495] = '{32'hc1843590, 32'hc1ffdba4, 32'hc2a5614d, 32'h40544745, 32'h41db025b, 32'h4232e4b9, 32'hc295acd7, 32'h428683ae};
test_label[4561] = '{32'hc2a5614d};
test_output[4561] = '{32'h4315f27e};
/*############ DEBUG ############
test_input[36488:36495] = '{-16.526153476, -31.9822462886, -82.6900410807, 3.3168498864, 27.3761509795, 44.7233631279, -74.8375775989, 67.2571892377};
test_label[4561] = '{-82.6900410807};
test_output[4561] = '{149.947230319};
############ END DEBUG ############*/
test_input[36496:36503] = '{32'h42a54f4c, 32'h42ba85aa, 32'hbfb22a73, 32'h4256cb4b, 32'h42c18e9c, 32'hc25956ad, 32'h4194c698, 32'hc22a1b5f};
test_label[4562] = '{32'h4256cb4b};
test_output[4562] = '{32'h422c6fde};
/*############ DEBUG ############
test_input[36496:36503] = '{82.6548770918, 93.2610593736, -1.39192045135, 53.6985300858, 96.7785309962, -54.3346459118, 18.59696883, -42.5267300049};
test_label[4562] = '{53.6985300858};
test_output[4562] = '{43.1092442291};
############ END DEBUG ############*/
test_input[36504:36511] = '{32'hc2758aea, 32'h42bdb89b, 32'h411f6779, 32'h42a05688, 32'hc2c70ffb, 32'hc2b95660, 32'hc1d53671, 32'hc28dfb99};
test_label[4563] = '{32'hc2b95660};
test_output[4563] = '{32'h433b877e};
/*############ DEBUG ############
test_input[36504:36511] = '{-61.3856564722, 94.8605578077, 9.96276175758, 80.1690054484, -99.5312146913, -92.6687025919, -26.6515825628, -70.9914000681};
test_label[4563] = '{-92.6687025919};
test_output[4563] = '{187.529260816};
############ END DEBUG ############*/
test_input[36512:36519] = '{32'hc24ac0d3, 32'hc20e355b, 32'hc24e6610, 32'hc2b7e13b, 32'h42aac1fd, 32'h42acfd24, 32'hc131aabb, 32'hc29e66a5};
test_label[4564] = '{32'hc2b7e13b};
test_output[4564] = '{32'h4332b7c2};
/*############ DEBUG ############
test_input[36512:36519] = '{-50.6883038323, -35.5521054245, -51.5996701887, -91.9399045531, 85.378880198, 86.4944131235, -11.1041823835, -79.200474163};
test_label[4564] = '{-91.9399045531};
test_output[4564] = '{178.717796355};
############ END DEBUG ############*/
test_input[36520:36527] = '{32'h41c163cc, 32'hc1c45f90, 32'h422f7828, 32'hc29ba2b3, 32'h419af8e7, 32'hc29bbb7b, 32'hc28302dc, 32'h4131c447};
test_label[4565] = '{32'h422f7828};
test_output[4565] = '{32'h3142006a};
/*############ DEBUG ############
test_input[36520:36527] = '{24.1737294483, -24.5466605282, 43.8673417466, -77.8177691039, 19.3715342147, -77.8661711208, -65.5055819178, 11.110419689};
test_label[4565] = '{43.8673417466};
test_output[4565] = '{2.82309498399e-09};
############ END DEBUG ############*/
test_input[36528:36535] = '{32'h42c17fe2, 32'hc2991f5c, 32'h4286befb, 32'hc1d4a90f, 32'hc20ebc62, 32'h41943bbc, 32'hc17cda69, 32'hc22c1995};
test_label[4566] = '{32'h41943bbc};
test_output[4566] = '{32'h429c70f3};
/*############ DEBUG ############
test_input[36528:36535] = '{96.749771802, -76.5612510215, 67.3730049306, -26.5825488013, -35.6839679258, 18.5291666901, -15.8033230776, -43.0249829303};
test_label[4566] = '{18.5291666901};
test_output[4566] = '{78.2206051119};
############ END DEBUG ############*/
test_input[36536:36543] = '{32'hc2c23f0a, 32'hc241b75e, 32'h41f4c3c9, 32'hc150c082, 32'hc2b3f4a7, 32'h41c14f6b, 32'h42b7cb25, 32'h42aeac4e};
test_label[4567] = '{32'hc2b3f4a7};
test_output[4567] = '{32'h4335e290};
/*############ DEBUG ############
test_input[36536:36543] = '{-97.1231264983, -48.4290699642, 30.5955973878, -13.0469990546, -89.9778353655, 24.1637791391, 91.8967641399, 87.3365339055};
test_label[4567] = '{-89.9778353655};
test_output[4567] = '{181.885004832};
############ END DEBUG ############*/
test_input[36544:36551] = '{32'hc22a3742, 32'hc19fe392, 32'hc0eeee39, 32'hc2c1e404, 32'h4199d4d8, 32'h415cd689, 32'h42993af4, 32'h40de4461};
test_label[4568] = '{32'hc0eeee39};
test_output[4568] = '{32'h42a829d7};
/*############ DEBUG ############
test_input[36544:36551] = '{-42.5539615614, -19.9861182376, -7.46657993339, -96.9453418615, 19.2289283995, 13.8023763825, 76.6151422344, 6.94584726208};
test_label[4568] = '{-7.46657993339};
test_output[4568] = '{84.0817221678};
############ END DEBUG ############*/
test_input[36552:36559] = '{32'h413fb010, 32'h429a0171, 32'h41f8ad5b, 32'hc2ad0d1c, 32'h401b0335, 32'h41a3a708, 32'hc1bddfa3, 32'h41aab5a2};
test_label[4569] = '{32'h401b0335};
test_output[4569] = '{32'h42952957};
/*############ DEBUG ############
test_input[36552:36559] = '{11.9804839594, 77.0028161932, 31.0846469732, -86.5256040413, 2.42207081692, 20.4565589673, -23.7341970185, 21.3386873449};
test_label[4569] = '{2.42207081692};
test_output[4569] = '{74.5807453763};
############ END DEBUG ############*/
test_input[36560:36567] = '{32'hc2b8d7c4, 32'h428cf0fe, 32'hc04081d4, 32'h4296b54c, 32'h41f65eac, 32'hc2312561, 32'hc25656eb, 32'h42b59d01};
test_label[4570] = '{32'h428cf0fe};
test_output[4570] = '{32'h41a2b00c};
/*############ DEBUG ############
test_input[36560:36567] = '{-92.4214148976, 70.4706888225, -3.00792404604, 75.354097643, 30.7962265569, -44.2865030874, -53.5848826183, 90.8066499007};
test_label[4570] = '{70.4706888225};
test_output[4570] = '{20.3359612742};
############ END DEBUG ############*/
test_input[36568:36575] = '{32'hc25e7056, 32'h42478a9d, 32'h42829e82, 32'hc27248e1, 32'h41a68909, 32'h42c006da, 32'hc22d26f9, 32'h425d95a1};
test_label[4571] = '{32'h41a68909};
test_output[4571] = '{32'h42966497};
/*############ DEBUG ############
test_input[36568:36575] = '{-55.609703282, 49.8853633785, 65.309582809, -60.5711726618, 20.816911029, 96.0133789827, -43.2880588513, 55.3961226537};
test_label[4571] = '{20.816911029};
test_output[4571] = '{75.1964679537};
############ END DEBUG ############*/
test_input[36576:36583] = '{32'h41a608f4, 32'h4202e7c8, 32'hc0f16d86, 32'hc249a6bb, 32'hc23a01b2, 32'hc299fc70, 32'h4211023a, 32'h428f7fdf};
test_label[4572] = '{32'hc299fc70};
test_output[4572] = '{32'h4314be28};
/*############ DEBUG ############
test_input[36576:36583] = '{20.7543711142, 32.7263504577, -7.54461943895, -50.4128230017, -46.5016557146, -76.9930450411, 36.2521750988, 71.7497511118};
test_label[4572] = '{-76.9930450411};
test_output[4572] = '{148.742796153};
############ END DEBUG ############*/
test_input[36584:36591] = '{32'hc28ad3b5, 32'h421538de, 32'h41936ab2, 32'hc10f0172, 32'h41aa70f9, 32'hc1e8f5a9, 32'hc263bda2, 32'hc2b537d8};
test_label[4573] = '{32'h41aa70f9};
test_output[4573] = '{32'h418000c2};
/*############ DEBUG ############
test_input[36584:36591] = '{-69.4134912699, 37.3055330756, 18.4270979437, -8.93785240345, 21.3051629346, -29.1199510065, -56.9351884614, -90.6090716723};
test_label[4573] = '{21.3051629346};
test_output[4573] = '{16.0003702597};
############ END DEBUG ############*/
test_input[36592:36599] = '{32'h41d5bd59, 32'h4286fbb4, 32'h418c7f6d, 32'h42936c4d, 32'hc271365b, 32'h4259744f, 32'hc2120e98, 32'hc2b7763a};
test_label[4574] = '{32'h42936c4d};
test_output[4574] = '{32'h3b023fc2};
/*############ DEBUG ############
test_input[36592:36599] = '{26.7174545318, 67.4916111516, 17.5622190173, 73.7115257098, -60.3030799072, 54.3635827184, -36.5142519583, -91.7309128904};
test_label[4574] = '{73.7115257098};
test_output[4574] = '{0.00198744287188};
############ END DEBUG ############*/
test_input[36600:36607] = '{32'hc2447b1f, 32'hc1dade7b, 32'h42b0b1b8, 32'hc23a0858, 32'h41a46e7d, 32'h42c7c618, 32'h42484a7f, 32'h426be303};
test_label[4575] = '{32'hc23a0858};
test_output[4575] = '{32'h43126522};
/*############ DEBUG ############
test_input[36600:36607] = '{-49.1202363796, -27.3586328783, 88.3471080337, -46.5081476633, 20.5539485553, 99.8869001194, 50.0727494354, 58.9716916757};
test_label[4575] = '{-46.5081476633};
test_output[4575] = '{146.395057517};
############ END DEBUG ############*/
test_input[36608:36615] = '{32'h41c055b4, 32'hc2638790, 32'h41b8f5a3, 32'h412fb44f, 32'hc21ed736, 32'h4280715d, 32'h42c1c75b, 32'hc2bf918d};
test_label[4576] = '{32'h41b8f5a3};
test_output[4576] = '{32'h429389f2};
/*############ DEBUG ############
test_input[36608:36615] = '{24.0418464326, -56.8823858665, 23.1199396772, 10.9815207048, -39.710167981, 64.2214090911, 96.8893628, -95.7842785161};
test_label[4576] = '{23.1199396772};
test_output[4576] = '{73.7694231228};
############ END DEBUG ############*/
test_input[36616:36623] = '{32'h42c22fb7, 32'hc23c6b50, 32'h41a3b5a1, 32'h429d3aa4, 32'h42495811, 32'hc20e0f32, 32'hc1afe43a, 32'hc2bafafd};
test_label[4577] = '{32'h42c22fb7};
test_output[4577] = '{32'h32221ee6};
/*############ DEBUG ############
test_input[36616:36623] = '{97.0931946146, -47.1047971361, 20.4636865043, 78.6145316032, 50.3360031139, -35.5148388592, -21.9864382404, -93.4902125232};
test_label[4577] = '{97.0931946146};
test_output[4577] = '{9.43666682585e-09};
############ END DEBUG ############*/
test_input[36624:36631] = '{32'h42788a31, 32'hc26bebdc, 32'h4239ffb9, 32'h4224e982, 32'h4290fcfa, 32'h42c1cbc6, 32'h423291cc, 32'hc285651f};
test_label[4578] = '{32'hc285651f};
test_output[4578] = '{32'h43239872};
/*############ DEBUG ############
test_input[36624:36631] = '{62.1349538569, -58.9803295737, 46.4997281181, 41.2280348528, 72.4940974231, 96.8979955442, 44.6423794407, -66.6975005297};
test_label[4578] = '{-66.6975005297};
test_output[4578] = '{163.595496074};
############ END DEBUG ############*/
test_input[36632:36639] = '{32'h42621ff2, 32'hc2a6fe09, 32'hc27d4ca5, 32'hc274f3ec, 32'hc1dd55f6, 32'hc2037a7c, 32'hc28e0aa8, 32'hc2a49389};
test_label[4579] = '{32'hc2a49389};
test_output[4579] = '{32'h430ad1c1};
/*############ DEBUG ############
test_input[36632:36639] = '{56.5311961485, -83.496163886, -63.3248484526, -61.2382062031, -27.6669735029, -32.8696122477, -71.0208137008, -82.2881518786};
test_label[4579] = '{-82.2881518786};
test_output[4579] = '{138.819348027};
############ END DEBUG ############*/
test_input[36640:36647] = '{32'hc2c450e3, 32'hc1a5070e, 32'hc235dd84, 32'h42006eca, 32'h42804584, 32'hc257547c, 32'hc262bf2f, 32'h42811296};
test_label[4580] = '{32'h42811296};
test_output[4580] = '{32'h3f034733};
/*############ DEBUG ############
test_input[36640:36647] = '{-98.1579801145, -20.6284439348, -45.4663240817, 32.1081941909, 64.1357741671, -53.8325027209, -56.6867038352, 64.5362978267};
test_label[4580] = '{64.5362978267};
test_output[4580] = '{0.512805134291};
############ END DEBUG ############*/
test_input[36648:36655] = '{32'hc08edd59, 32'h41e9333d, 32'hc2b262b1, 32'h41f93b6e, 32'h41148808, 32'hc1b902cf, 32'h413ec9c9, 32'hc2aa16ee};
test_label[4581] = '{32'h413ec9c9};
test_output[4581] = '{32'h419ad983};
/*############ DEBUG ############
test_input[36648:36655] = '{-4.46451995881, 29.1500192325, -89.1927588666, 31.1540187414, 9.28321078074, -23.1263704948, 11.9242640029, -85.0447882928};
test_label[4581] = '{11.9242640029};
test_output[4581] = '{19.3562068395};
############ END DEBUG ############*/
test_input[36656:36663] = '{32'hc1e901b6, 32'hc28129d9, 32'h42a164ea, 32'h429c69ac, 32'h4138e9d0, 32'hc211323d, 32'h42c186b2, 32'hc009def5};
test_label[4582] = '{32'h42a164ea};
test_output[4582] = '{32'h41808720};
/*############ DEBUG ############
test_input[36656:36663] = '{-29.1258352417, -64.5817332017, 80.6971002334, 78.2063900205, 11.5570834519, -36.2990609253, 96.7630796527, -2.15423331309};
test_label[4582] = '{80.6971002334};
test_output[4582] = '{16.0659795334};
############ END DEBUG ############*/
test_input[36664:36671] = '{32'hc2505c53, 32'hc05f45b7, 32'h422e11ff, 32'hc20bfa5b, 32'hc19f1ad8, 32'h423cf10d, 32'h42870888, 32'h4291b975};
test_label[4583] = '{32'hc05f45b7};
test_output[4583] = '{32'h4298b612};
/*############ DEBUG ############
test_input[36664:36671] = '{-52.0901590102, -3.48863007746, 43.5175737295, -34.9944866808, -19.8881067873, 47.2354011154, 67.5166603174, 72.8622211177};
test_label[4583] = '{-3.48863007746};
test_output[4583] = '{76.3556091341};
############ END DEBUG ############*/
test_input[36672:36679] = '{32'h428154e6, 32'hc1eb8652, 32'hc23f6e0c, 32'h42082158, 32'h41f815c1, 32'h41184ea3, 32'h41804082, 32'hc2a240eb};
test_label[4584] = '{32'hc1eb8652};
test_output[4584] = '{32'h42bc367b};
/*############ DEBUG ############
test_input[36672:36679] = '{64.6658183912, -29.4405865775, -47.8574672224, 34.0325636954, 31.0106217253, 9.51919888385, 16.0314984434, -81.1267909014};
test_label[4584] = '{-29.4405865775};
test_output[4584] = '{94.1064049687};
############ END DEBUG ############*/
test_input[36680:36687] = '{32'hc1d5ffc8, 32'h4267fb26, 32'hc2aac2d4, 32'hc27705cc, 32'h42bc3e81, 32'h3fa5b1e0, 32'hc22449af, 32'h42940c01};
test_label[4585] = '{32'hc22449af};
test_output[4585] = '{32'h430731ac};
/*############ DEBUG ############
test_input[36680:36687] = '{-26.7498934214, 57.9952624069, -85.3805251792, -61.7556619587, 94.1220787823, 1.29449075493, -41.0719559726, 74.0234465808};
test_label[4585] = '{-41.0719559726};
test_output[4585] = '{135.194034757};
############ END DEBUG ############*/
test_input[36688:36695] = '{32'h42517600, 32'h42a6a0ff, 32'h41c346aa, 32'hc1b12cdf, 32'h420fe316, 32'hc1f26847, 32'h42b12eb8, 32'h42b112e8};
test_label[4586] = '{32'h41c346aa};
test_output[4586] = '{32'h4281b391};
/*############ DEBUG ############
test_input[36688:36695] = '{52.3652327552, 83.3144457037, 24.4095040163, -22.146909743, 35.9717631055, -30.3009174625, 88.5912448782, 88.5369269446};
test_label[4586] = '{24.4095040163};
test_output[4586] = '{64.8507181347};
############ END DEBUG ############*/
test_input[36696:36703] = '{32'h42b37a8b, 32'h42295fbe, 32'h42a8a1fb, 32'h4288b4bc, 32'h42bdf1a0, 32'h42b393e1, 32'hc1a662c0, 32'h41f03cb1};
test_label[4587] = '{32'h42b37a8b};
test_output[4587] = '{32'h40a7cab5};
/*############ DEBUG ############
test_input[36696:36703] = '{89.7393409393, 42.3434991072, 84.3163643087, 68.3530000628, 94.9719211753, 89.7888256184, -20.7982173305, 30.0296347828};
test_label[4587] = '{89.7393409393};
test_output[4587] = '{5.24349437038};
############ END DEBUG ############*/
test_input[36704:36711] = '{32'h42c34dbe, 32'h41b02a26, 32'h421fb120, 32'h42adc58e, 32'h42c64c2d, 32'h42213f49, 32'h410c49f9, 32'hc2b884bb};
test_label[4588] = '{32'h41b02a26};
test_output[4588] = '{32'h429aa90d};
/*############ DEBUG ############
test_input[36704:36711] = '{97.6518364677, 22.0205807331, 39.9229741937, 86.8858527684, 99.1487818147, 40.3118026024, 8.76805959683, -92.2592382032};
test_label[4588] = '{22.0205807331};
test_output[4588] = '{77.3301761623};
############ END DEBUG ############*/
test_input[36712:36719] = '{32'hc2b64c82, 32'h41592018, 32'hc29f00a1, 32'hc21a5c0c, 32'hc1c92bf9, 32'h42aaae77, 32'hc03e841a, 32'h424889fa};
test_label[4589] = '{32'hc2b64c82};
test_output[4589] = '{32'h43307d7c};
/*############ DEBUG ############
test_input[36712:36719] = '{-91.1494255703, 13.5703358158, -79.5012280973, -38.5898887285, -25.1464702089, 85.3407550976, -2.97681284479, 50.1347410542};
test_label[4589] = '{-91.1494255703};
test_output[4589] = '{176.490180668};
############ END DEBUG ############*/
test_input[36720:36727] = '{32'hc1c94fc2, 32'h429af2f0, 32'hc2af8a01, 32'h4188b8e8, 32'h427fb564, 32'hc1212eed, 32'hc131a422, 32'hc0e0baba};
test_label[4590] = '{32'hc131a422};
test_output[4590] = '{32'h42b12774};
/*############ DEBUG ############
test_input[36720:36727] = '{-25.1639441825, 77.4744848453, -87.7695351371, 17.0902860689, 63.9271399509, -10.0739567509, -11.1025711082, -7.0227935634};
test_label[4590] = '{-11.1025711082};
test_output[4590] = '{88.5770572611};
############ END DEBUG ############*/
test_input[36728:36735] = '{32'h429fee18, 32'hc22f9b49, 32'h4043a379, 32'hc2bb399d, 32'hc2015c8e, 32'h42368e18, 32'hc2443c87, 32'h41b795fb};
test_label[4591] = '{32'hc2bb399d};
test_output[4591] = '{32'h432d93da};
/*############ DEBUG ############
test_input[36728:36735] = '{79.9650247153, -43.9016451642, 3.0568526337, -93.6125237087, -32.3403836249, 45.6387618306, -49.0591081947, 22.9482324309};
test_label[4591] = '{-93.6125237087};
test_output[4591] = '{173.577548424};
############ END DEBUG ############*/
test_input[36736:36743] = '{32'h42ba83d1, 32'hc1b55b6a, 32'h42254e01, 32'h4208923b, 32'hc26923a8, 32'hc22a381a, 32'hc18b702f, 32'h42c7080a};
test_label[4592] = '{32'h4208923b};
test_output[4592] = '{32'h4282bfe7};
/*############ DEBUG ############
test_input[36736:36743] = '{93.2574543491, -22.6696360203, 41.3261756878, 34.1428050591, -58.2848190553, -42.5547862589, -17.4297762631, 99.5157041968};
test_label[4592] = '{34.1428050591};
test_output[4592] = '{65.374811901};
############ END DEBUG ############*/
test_input[36744:36751] = '{32'h420811ab, 32'hc282ae50, 32'h402e441a, 32'hc04a2405, 32'h425855ac, 32'hc0fcc3cd, 32'hc2035147, 32'h42c716bc};
test_label[4593] = '{32'h420811ab};
test_output[4593] = '{32'h42830de7};
/*############ DEBUG ############
test_input[36744:36751] = '{34.0172546752, -65.3404547466, 2.7229066965, -3.15844837314, 54.0836639339, -7.898901245, -32.8293713558, 99.5444047198};
test_label[4593] = '{34.0172546752};
test_output[4593] = '{65.5271500445};
############ END DEBUG ############*/
test_input[36752:36759] = '{32'hc1add021, 32'hc13197d2, 32'hc28586d9, 32'hc0dbefd1, 32'hc25f0e68, 32'h4093d141, 32'hc2072f04, 32'hc2036ed3};
test_label[4594] = '{32'hc28586d9};
test_output[4594] = '{32'h428ec3ef};
/*############ DEBUG ############
test_input[36752:36759] = '{-21.7266258375, -11.0995653053, -66.7633749327, -6.8730245388, -55.7640704613, 4.61929390714, -33.7959131281, -32.8582256439};
test_label[4594] = '{-66.7633749327};
test_output[4594] = '{71.3826791971};
############ END DEBUG ############*/
test_input[36760:36767] = '{32'hc1da462b, 32'hc25d411b, 32'h429284f3, 32'h41d50609, 32'hc299f1b0, 32'hc2a581ff, 32'h4146cbda, 32'h4137f79a};
test_label[4595] = '{32'hc299f1b0};
test_output[4595] = '{32'h43163b51};
/*############ DEBUG ############
test_input[36760:36767] = '{-27.2842610107, -55.3135811403, 73.2596645359, 26.6279475755, -76.9720447253, -82.7538963936, 12.4247679928, 11.4979493034};
test_label[4595] = '{-76.9720447253};
test_output[4595] = '{150.231709261};
############ END DEBUG ############*/
test_input[36768:36775] = '{32'h416bb015, 32'h426b1673, 32'hc2a15d3c, 32'h425eaa59, 32'hc1fd4c46, 32'h4228a7c6, 32'h42ab9b52, 32'hc21275c3};
test_label[4596] = '{32'hc1fd4c46};
test_output[4596] = '{32'h42eaee63};
/*############ DEBUG ############
test_input[36768:36775] = '{14.7304885522, 58.7719245096, -80.6820981271, 55.6663559791, -31.6622424319, 42.1638402088, 85.8033601413, -36.6150034906};
test_label[4596] = '{-31.6622424319};
test_output[4596] = '{117.465602573};
############ END DEBUG ############*/
test_input[36776:36783] = '{32'h427987d3, 32'h41a9705b, 32'h41eeb37b, 32'hc2c154f1, 32'hc2c003fb, 32'hc0b47897, 32'hc1f0beb1, 32'h42c27122};
test_label[4597] = '{32'hc1f0beb1};
test_output[4597] = '{32'h42fea0ce};
/*############ DEBUG ############
test_input[36776:36783] = '{62.3826404906, 21.1798602675, 29.837636427, -96.6658993773, -96.0077769162, -5.63972044531, -30.0931109115, 97.220963112};
test_label[4597] = '{-30.0931109115};
test_output[4597] = '{127.314074024};
############ END DEBUG ############*/
test_input[36784:36791] = '{32'hc0da37ac, 32'hc2bbf4bd, 32'hc2163bcd, 32'hc1adc1df, 32'hc2b6be5c, 32'h42359fa2, 32'hc1935065, 32'hc27c832d};
test_label[4598] = '{32'hc0da37ac};
test_output[4598] = '{32'h4250e697};
/*############ DEBUG ############
test_input[36784:36791] = '{-6.81929576062, -93.9780066892, -37.5583986763, -21.7196630039, -91.3717944288, 45.405891528, -18.4142554671, -63.1281002075};
test_label[4598] = '{-6.81929576062};
test_output[4598] = '{52.2251872886};
############ END DEBUG ############*/
test_input[36792:36799] = '{32'hc24f13d7, 32'h4094a45b, 32'hc227a1b0, 32'h41984794, 32'hc005811a, 32'h42a0a79d, 32'hc299bcf7, 32'hc20b61e1};
test_label[4599] = '{32'h42a0a79d};
test_output[4599] = '{32'h80000000};
/*############ DEBUG ############
test_input[36792:36799] = '{-51.7693743639, 4.64506307891, -41.907898322, 19.0349494708, -2.08600485139, 80.327372887, -76.8690698487, -34.8455843212};
test_label[4599] = '{80.327372887};
test_output[4599] = '{-0.0};
############ END DEBUG ############*/
test_input[36800:36807] = '{32'h420ca7b6, 32'h41db3df0, 32'h41930ab2, 32'hc2ac8b09, 32'h401e0d93, 32'hc278880f, 32'h42189d9a, 32'hc2af220a};
test_label[4600] = '{32'hc2af220a};
test_output[4600] = '{32'h42fb89f7};
/*############ DEBUG ############
test_input[36800:36807] = '{35.1637808688, 27.4052436399, 18.3802232477, -86.2715556017, 2.46957849371, -62.132869843, 38.1539065558, -87.5664787608};
test_label[4600] = '{-87.5664787608};
test_output[4600] = '{125.769463623};
############ END DEBUG ############*/
test_input[36808:36815] = '{32'h42a4ba13, 32'hc264f9c1, 32'hc239f23f, 32'h42ba2a6d, 32'h42a92801, 32'hc292735f, 32'h417a750f, 32'hc1cd798b};
test_label[4601] = '{32'hc239f23f};
test_output[4601] = '{32'h430b91d5};
/*############ DEBUG ############
test_input[36808:36815] = '{82.3634247672, -57.2439002027, -46.4865679873, 93.082863641, 84.578135269, -73.2253372026, 15.6535790462, -25.6843462798};
test_label[4601] = '{-46.4865679873};
test_output[4601] = '{139.569656223};
############ END DEBUG ############*/
test_input[36816:36823] = '{32'h4126a770, 32'h4287e001, 32'hc29777ed, 32'hc06e93ef, 32'h42838dd5, 32'h42c5715b, 32'hc2b74552, 32'h4284f197};
test_label[4602] = '{32'h42c5715b};
test_output[4602] = '{32'h29818000};
/*############ DEBUG ############
test_input[36816:36823] = '{10.4158782529, 67.937507428, -75.7342263976, -3.72777920795, 65.7770140611, 98.721400963, -91.6353881988, 66.4718584413};
test_label[4602] = '{98.721400963};
test_output[4602] = '{5.75095526756e-14};
############ END DEBUG ############*/
test_input[36824:36831] = '{32'h42b8cf80, 32'h4289a4e3, 32'h41d313e3, 32'h404f97c2, 32'hc2b6578e, 32'h4228771a, 32'hc25e0c25, 32'hc2a96a32};
test_label[4603] = '{32'h404f97c2};
test_output[4603] = '{32'h42b252c2};
/*############ DEBUG ############
test_input[36824:36831] = '{92.4052721173, 68.8220407551, 26.3847108321, 3.24363748288, -91.1710064213, 42.1163086895, -55.5118608166, -84.707411527};
test_label[4603] = '{3.24363748288};
test_output[4603] = '{89.1616346345};
############ END DEBUG ############*/
test_input[36832:36839] = '{32'hc189cbc5, 32'h420b03fa, 32'h42064dcd, 32'h41c10ec6, 32'h428ca8bb, 32'hc196b19b, 32'h3f4bacc8, 32'hc2afe543};
test_label[4604] = '{32'hc196b19b};
test_output[4604] = '{32'h42b25521};
/*############ DEBUG ############
test_input[36832:36839] = '{-17.224496064, 34.7538849069, 33.575978055, 24.1322132595, 70.3295487285, -18.8367217424, 0.79560516036, -87.9477778271};
test_label[4604] = '{-18.8367217424};
test_output[4604] = '{89.1662704709};
############ END DEBUG ############*/
test_input[36840:36847] = '{32'hc1ddbf54, 32'hc0a4fb6f, 32'h42802283, 32'h4174f46a, 32'h3f13764c, 32'h42a23634, 32'h4196f33e, 32'hc29fbdc4};
test_label[4605] = '{32'h3f13764c};
test_output[4605] = '{32'h42a10f47};
/*############ DEBUG ############
test_input[36840:36847] = '{-27.7184221296, -5.15569248349, 64.0674085652, 15.3096711017, 0.576023817236, 81.1058655201, 18.8687709531, -79.8706349678};
test_label[4605] = '{0.576023817236};
test_output[4605] = '{80.5298417427};
############ END DEBUG ############*/
test_input[36848:36855] = '{32'hc25b03fa, 32'h424a1b7c, 32'hc28bb008, 32'h428053d3, 32'h42a535f2, 32'hc2926353, 32'hc074770d, 32'hc299511c};
test_label[4606] = '{32'hc25b03fa};
test_output[4606] = '{32'h43095bf7};
/*############ DEBUG ############
test_input[36848:36855] = '{-54.7538847153, 50.5268402673, -69.8438090248, 64.1637213912, 82.6053597119, -73.1939917865, -3.81976631512, -76.6584130513};
test_label[4606] = '{-54.7538847153};
test_output[4606] = '{137.359244437};
############ END DEBUG ############*/
test_input[36856:36863] = '{32'h42b53a74, 32'h42993e41, 32'hc2702b68, 32'hc1ec9f17, 32'h429a5e75, 32'h423886a5, 32'h409f5c38, 32'h42c2afb2};
test_label[4607] = '{32'hc2702b68};
test_output[4607] = '{32'h431d6301};
/*############ DEBUG ############
test_input[36856:36863] = '{90.6141663277, 76.6215858612, -60.0423874658, -29.5776797137, 77.1844895358, 46.1314888618, 4.98000698383, 97.3431574469};
test_label[4607] = '{-60.0423874658};
test_output[4607] = '{157.38673994};
############ END DEBUG ############*/
test_input[36864:36871] = '{32'hc27745b2, 32'h4006fe70, 32'h4228b2a2, 32'h4291db69, 32'hc26ad9c8, 32'hc1f6f6b0, 32'h42c0ae46, 32'hc293b4c6};
test_label[4608] = '{32'hc293b4c6};
test_output[4608] = '{32'h432a3186};
/*############ DEBUG ############
test_input[36864:36871] = '{-61.8180603684, 2.10927957734, 42.174445429, 72.9285382019, -58.7126766384, -30.8704532564, 96.3403774692, -73.8530714888};
test_label[4608] = '{-73.8530714888};
test_output[4608] = '{170.193448958};
############ END DEBUG ############*/
test_input[36872:36879] = '{32'h413a2c5e, 32'h418f5b7c, 32'h42ac229d, 32'hc0dc3239, 32'h42ab3695, 32'h42b83796, 32'hc2431d82, 32'h42bb0a22};
test_label[4609] = '{32'h418f5b7c};
test_output[4609] = '{32'h4297a35f};
/*############ DEBUG ############
test_input[36872:36879] = '{11.6358313802, 17.9196699419, 86.0676073597, -6.88113046871, 85.6066071202, 92.1085649919, -48.7788180223, 93.5197902993};
test_label[4609] = '{17.9196699419};
test_output[4609] = '{75.8190875017};
############ END DEBUG ############*/
test_input[36880:36887] = '{32'hc27c8999, 32'hc2b3035d, 32'hc27f7489, 32'hc0ca831c, 32'hc2b15333, 32'hc225a046, 32'hc280d85c, 32'hc19ca1e9};
test_label[4610] = '{32'hc27f7489};
test_output[4610] = '{32'h42662426};
/*############ DEBUG ############
test_input[36880:36887] = '{-63.1343723511, -89.5065668109, -63.8638037155, -6.32850445878, -88.6624952131, -41.4065162405, -64.4225788624, -19.5790578415};
test_label[4610] = '{-63.8638037155};
test_output[4610] = '{57.5353010161};
############ END DEBUG ############*/
test_input[36888:36895] = '{32'hc28de2e3, 32'hc2c368c6, 32'h42502084, 32'hc20b8aa0, 32'h3f8d7876, 32'h413720e3, 32'hc2a07468, 32'hc2a01720};
test_label[4611] = '{32'h3f8d7876};
test_output[4611] = '{32'h424bb4c0};
/*############ DEBUG ############
test_input[36888:36895] = '{-70.9431396567, -97.7046384278, 52.0317517141, -34.8853778447, 1.10523868033, 11.4455289434, -80.227358343, -80.0451697079};
test_label[4611] = '{1.10523868033};
test_output[4611] = '{50.9265130337};
############ END DEBUG ############*/
test_input[36896:36903] = '{32'hc2a0c1dd, 32'hc27e7eeb, 32'h419d9e84, 32'h420f7559, 32'hc1314e61, 32'hc18d480b, 32'h4291914a, 32'hc2a321fa};
test_label[4612] = '{32'h420f7559};
test_output[4612] = '{32'h4213ad3b};
/*############ DEBUG ############
test_input[36896:36903] = '{-80.3786388783, -63.6239417838, 19.7024005131, 35.864598095, -11.0816352782, -17.660177733, 72.7837672203, -81.5663631864};
test_label[4612] = '{35.864598095};
test_output[4612] = '{36.9191691253};
############ END DEBUG ############*/
test_input[36904:36911] = '{32'h4289bcf9, 32'hc29bc4d7, 32'hc2716103, 32'hc2a8fbfc, 32'h414742ce, 32'hc281e13f, 32'h42b22471, 32'h42b2d86d};
test_label[4613] = '{32'h4289bcf9};
test_output[4613] = '{32'h41a8b0e2};
/*############ DEBUG ############
test_input[36904:36911] = '{68.8690895224, -77.8844521947, -60.3447389406, -84.4921541669, 12.4538096865, -64.939933593, 89.0711754691, 89.4227094271};
test_label[4613] = '{68.8690895224};
test_output[4613] = '{21.0863682348};
############ END DEBUG ############*/
test_input[36912:36919] = '{32'h408593ae, 32'h4240ce35, 32'h42064e34, 32'h421d2482, 32'hc248613e, 32'h4299be1f, 32'hc28a9245, 32'h428211c9};
test_label[4614] = '{32'h428211c9};
test_output[4614] = '{32'h413d62ba};
/*############ DEBUG ############
test_input[36912:36919] = '{4.17427712088, 48.2013736719, 33.5763687185, 39.2856515862, -50.0949619585, 76.8713305718, -69.2856831445, 65.0347348953};
test_label[4614] = '{65.0347348953};
test_output[4614] = '{11.8366029113};
############ END DEBUG ############*/
test_input[36920:36927] = '{32'hc207bc01, 32'hc1c9d1e5, 32'hc229b5ff, 32'h422d021f, 32'h427d02e1, 32'hc15df8c7, 32'hc25512bb, 32'h4206cdda};
test_label[4615] = '{32'hc207bc01};
test_output[4615] = '{32'h42c25f71};
/*############ DEBUG ############
test_input[36920:36927] = '{-33.9335985734, -25.2274868017, -42.4277300046, 43.2520700068, 63.252812143, -13.8732365806, -53.2682907056, 33.7010279691};
test_label[4615] = '{-33.9335985734};
test_output[4615] = '{97.1864107184};
############ END DEBUG ############*/
test_input[36928:36935] = '{32'h4298f6fd, 32'hc252390b, 32'h40e1fe24, 32'hc1de76c6, 32'hc2bb8f2b, 32'hc1d4d80f, 32'hc26c98c4, 32'h42bf11d3};
test_label[4616] = '{32'hc26c98c4};
test_output[4616] = '{32'h431aaf1a};
/*############ DEBUG ############
test_input[36928:36935] = '{76.4823963864, -52.5557063571, 7.06227299372, -27.8079950361, -93.7796252471, -26.6054966163, -59.149185672, 95.5348110065};
test_label[4616] = '{-59.149185672};
test_output[4616] = '{154.683996684};
############ END DEBUG ############*/
test_input[36936:36943] = '{32'hc1a3d785, 32'hc26302f7, 32'h4293dd20, 32'h421534fa, 32'h4284e642, 32'h42b5a6b6, 32'h409d0980, 32'hc20db1b2};
test_label[4617] = '{32'h421534fa};
test_output[4617] = '{32'h42561872};
/*############ DEBUG ############
test_input[36936:36943] = '{-20.4802337389, -56.7528969804, 73.931882181, 37.3017339669, 66.4497249623, 90.8256066177, 4.90740976296, -35.4235310361};
test_label[4617] = '{37.3017339669};
test_output[4617] = '{53.5238726968};
############ END DEBUG ############*/
test_input[36944:36951] = '{32'hc1e697ba, 32'hc2badfc8, 32'hc29229e5, 32'h42a5d5de, 32'hc16d9c1a, 32'hc2617b9c, 32'hc10c5f62, 32'h42a3e8ae};
test_label[4618] = '{32'hc2badfc8};
test_output[4618] = '{32'h4330ad95};
/*############ DEBUG ############
test_input[36944:36951] = '{-28.8240860764, -93.4370720035, -73.0818237287, 82.9177113807, -14.8506108901, -56.3707108546, -8.77328639081, 81.9544522396};
test_label[4618] = '{-93.4370720035};
test_output[4618] = '{176.678059661};
############ END DEBUG ############*/
test_input[36952:36959] = '{32'h42c295c4, 32'hc264c45c, 32'h4200c013, 32'h4231f406, 32'h420e6da8, 32'hc25f52c1, 32'h41b1a978, 32'h41875bb3};
test_label[4619] = '{32'h420e6da8};
test_output[4619] = '{32'h4276bde1};
/*############ DEBUG ############
test_input[36952:36959] = '{97.2925146035, -57.1917572196, 32.1875736892, 44.4883044599, 35.6070858529, -55.8308162613, 22.2077480986, 16.919775415};
test_label[4619] = '{35.6070858529};
test_output[4619] = '{61.6854287506};
############ END DEBUG ############*/
test_input[36960:36967] = '{32'h41a2e991, 32'h41f6c37a, 32'hc29529f3, 32'hc1e421e7, 32'hc29c6807, 32'h42a5242f, 32'hc2c768be, 32'hc1acaabb};
test_label[4620] = '{32'h42a5242f};
test_output[4620] = '{32'h80000000};
/*############ DEBUG ############
test_input[36960:36967] = '{20.3640469399, 30.845447884, -74.5819322712, -28.5165531612, -78.2031747945, 82.5706700798, -99.7045718085, -21.5833645777};
test_label[4620] = '{82.5706700798};
test_output[4620] = '{-0.0};
############ END DEBUG ############*/
test_input[36968:36975] = '{32'h4252566d, 32'hc2abf633, 32'hc1fee920, 32'h42a589c4, 32'h421548f2, 32'hc2870753, 32'hbf33ee03, 32'hc28dfbfe};
test_label[4621] = '{32'hc28dfbfe};
test_output[4621] = '{32'h4319c2e1};
/*############ DEBUG ############
test_input[36968:36975] = '{52.5844010841, -85.9808594895, -31.8638314905, 82.7690705893, 37.3212362888, -67.5143030965, -0.702850502381, -70.9921740432};
test_label[4621] = '{-70.9921740432};
test_output[4621] = '{153.761244632};
############ END DEBUG ############*/
test_input[36976:36983] = '{32'hc2a0487e, 32'h42960ec0, 32'hc25b9b86, 32'hc1425379, 32'hc14702cd, 32'h428058b3, 32'hc2c6d371, 32'hc2ab1c63};
test_label[4622] = '{32'hc2a0487e};
test_output[4622] = '{32'h431b2ba0};
/*############ DEBUG ############
test_input[36976:36983] = '{-80.1415849134, 75.0288080117, -54.9018778276, -12.1453788203, -12.438183979, 64.1732437784, -99.4129747315, -85.5554446714};
test_label[4622] = '{-80.1415849134};
test_output[4622] = '{155.170412222};
############ END DEBUG ############*/
test_input[36984:36991] = '{32'hc085fcfe, 32'hc098908c, 32'h42c5553e, 32'hc0ddac27, 32'hc2be85a5, 32'h42495098, 32'h42764601, 32'h42338f52};
test_label[4623] = '{32'hc2be85a5};
test_output[4623] = '{32'h4341ed71};
/*############ DEBUG ############
test_input[36984:36991] = '{-4.18713304033, -4.76764493024, 98.6664863032, -6.92726463502, -95.2610249683, 50.3287032041, 61.5683636589, 44.8899610239};
test_label[4623] = '{-95.2610249683};
test_output[4623] = '{193.927511272};
############ END DEBUG ############*/
test_input[36992:36999] = '{32'h41c22535, 32'h4106515a, 32'h41698891, 32'hc1c07616, 32'hc21881a0, 32'hc2a3c5d4, 32'h41ab4d30, 32'hc28c8da9};
test_label[4624] = '{32'hc1c07616};
test_output[4624] = '{32'h424186fc};
/*############ DEBUG ############
test_input[36992:36999] = '{24.268166769, 8.39486157095, 14.5958410255, -24.0576595335, -38.1265881746, -81.8863816313, 21.4126883823, -70.2766828713};
test_label[4624] = '{-24.0576595335};
test_output[4624] = '{48.3818203842};
############ END DEBUG ############*/
test_input[37000:37007] = '{32'h41809339, 32'hc2b328e6, 32'h42ac1c6d, 32'h426ca581, 32'h4284456e, 32'hc219f846, 32'hc2c63e13, 32'h4268400c};
test_label[4625] = '{32'h41809339};
test_output[4625] = '{32'h428bf79e};
/*############ DEBUG ############
test_input[37000:37007] = '{16.0718862503, -89.579882156, 86.055516087, 59.161625749, 66.1356061801, -38.4924544502, -99.1212378773, 58.0625442916};
test_label[4625] = '{16.0718862503};
test_output[4625] = '{69.9836298389};
############ END DEBUG ############*/
test_input[37008:37015] = '{32'h42a18e2e, 32'h42bf4f39, 32'h4289dd62, 32'hc29348f8, 32'hc29cb802, 32'hc265c95c, 32'h42a3540d, 32'hc22d2738};
test_label[4626] = '{32'hc22d2738};
test_output[4626] = '{32'h430af16a};
/*############ DEBUG ############
test_input[37008:37015] = '{80.7776915274, 95.6547300483, 68.9323911352, -73.6425143594, -78.3593922845, -57.4466399232, 81.6641647111, -43.2882987374};
test_label[4626] = '{-43.2882987374};
test_output[4626] = '{138.943029971};
############ END DEBUG ############*/
test_input[37016:37023] = '{32'hc1b75721, 32'hc2ad49a6, 32'hc28f2c67, 32'hc28b8810, 32'h3f0e22fd, 32'hc28e35ce, 32'h42aada75, 32'hc23d9ca0};
test_label[4627] = '{32'h3f0e22fd};
test_output[4627] = '{32'h42a9be2f};
/*############ DEBUG ############
test_input[37016:37023] = '{-22.9175426182, -86.6438436407, -71.5867208, -69.7657463669, 0.555221394874, -71.1050870587, 85.426676668, -47.4029537247};
test_label[4627] = '{0.555221394874};
test_output[4627] = '{84.8714552731};
############ END DEBUG ############*/
test_input[37024:37031] = '{32'hc2beae58, 32'hc2283d73, 32'h41aec05f, 32'hc1cd52cf, 32'h422faa4a, 32'hc161c344, 32'hc19cbe04, 32'hc02796a3};
test_label[4628] = '{32'hc19cbe04};
test_output[4628] = '{32'h427e094c};
/*############ DEBUG ############
test_input[37024:37031] = '{-95.3405185564, -42.0600078702, 21.8439320875, -25.6654334071, 43.9162966684, -14.1101722343, -19.5927813569, -2.61856916061};
test_label[4628] = '{-19.5927813569};
test_output[4628] = '{63.5090780256};
############ END DEBUG ############*/
test_input[37032:37039] = '{32'hc299c849, 32'h40c9a58e, 32'h429cabf2, 32'hc18bdc43, 32'hc065d409, 32'hc167dabc, 32'h41d3439e, 32'h42a0407d};
test_label[4629] = '{32'h41d3439e};
test_output[4629] = '{32'h42577d43};
/*############ DEBUG ############
test_input[37032:37039] = '{-76.8911854013, 6.30145950792, 78.3358342401, -17.4825499856, -3.59106667527, -14.4909016963, 26.408015319, 80.1259564088};
test_label[4629] = '{26.408015319};
test_output[4629] = '{53.8723258339};
############ END DEBUG ############*/
test_input[37040:37047] = '{32'h424f5b6d, 32'h42b6faf2, 32'h415b12c1, 32'h42475b82, 32'h41f246e4, 32'hc2bff767, 32'h42c6a436, 32'h41359601};
test_label[4630] = '{32'h415b12c1};
test_output[4630] = '{32'h42ab4212};
/*############ DEBUG ############
test_input[37040:37047] = '{51.8392814648, 91.4901281975, 13.6920788233, 49.8393626287, 30.2846137242, -95.9832098733, 99.320721717, 11.3491223382};
test_label[4630] = '{13.6920788233};
test_output[4630] = '{85.6290402044};
############ END DEBUG ############*/
test_input[37048:37055] = '{32'h41c24573, 32'hc2b230d7, 32'hc26e80fb, 32'hc1fa007b, 32'hc1943aba, 32'hbfe5d6a1, 32'h42c34f01, 32'h426bb2d1};
test_label[4631] = '{32'hc26e80fb};
test_output[4631] = '{32'h431d47bf};
/*############ DEBUG ############
test_input[37048:37055] = '{24.2839113085, -89.0953916002, -59.6259585565, -31.2502337329, -18.5286759076, -1.79561242198, 97.6543061311, 58.9246245905};
test_label[4631] = '{-59.6259585565};
test_output[4631] = '{157.280264688};
############ END DEBUG ############*/
test_input[37056:37063] = '{32'hc2be44ce, 32'h428020c6, 32'h41fa9876, 32'hc1fffd28, 32'hc25a1832, 32'h4270b164, 32'hc23a3fab, 32'hc01ba809};
test_label[4632] = '{32'hc23a3fab};
test_output[4632] = '{32'h42dd4af6};
/*############ DEBUG ############
test_input[37056:37063] = '{-95.1343805672, 64.0640091157, 31.324443027, -31.9986119625, -54.5236270062, 60.1732331344, -46.5621749099, -2.43213103776};
test_label[4632] = '{-46.5621749099};
test_output[4632] = '{110.64640763};
############ END DEBUG ############*/
test_input[37064:37071] = '{32'hc2a8f9b3, 32'h421ba8b2, 32'hc1bd84a5, 32'hc2a9d792, 32'h42575a33, 32'hc08a7895, 32'hc2379a7d, 32'hc2046945};
test_label[4633] = '{32'hc1bd84a5};
test_output[4633] = '{32'h429b0e43};
/*############ DEBUG ############
test_input[37064:37071] = '{-84.4876913726, 38.9147416366, -23.6897685387, -84.9210353441, 53.838086213, -4.32721950916, -45.9008683933, -33.1028008718};
test_label[4633] = '{-23.6897685387};
test_output[4633] = '{77.5278550819};
############ END DEBUG ############*/
test_input[37072:37079] = '{32'h42a50c78, 32'hc29f1ed0, 32'hc2b62f18, 32'h42072f85, 32'h420bf256, 32'h40b1367c, 32'h4266f739, 32'hc240661b};
test_label[4634] = '{32'h420bf256};
test_output[4634] = '{32'h423e269a};
/*############ DEBUG ############
test_input[37072:37079] = '{82.5243538418, -79.5601822791, -91.0919816829, 33.7964061979, 34.9866575362, 5.53790090029, 57.7414292402, -48.0997142314};
test_label[4634] = '{34.9866575362};
test_output[4634] = '{47.5376963056};
############ END DEBUG ############*/
test_input[37080:37087] = '{32'hc067e405, 32'hc2bca880, 32'h400bdd54, 32'h4265458a, 32'h41b39461, 32'hc2953243, 32'h42a9cb4e, 32'hbebb9e37};
test_label[4635] = '{32'h41b39461};
test_output[4635] = '{32'h4279cc6c};
/*############ DEBUG ############
test_input[37080:37087] = '{-3.62329215166, -94.3291019224, 2.18538382587, 57.3179083513, 22.4474504502, -74.5981689678, 84.8970797724, -0.36644144677};
test_label[4635] = '{22.4474504502};
test_output[4635] = '{62.4496293222};
############ END DEBUG ############*/
test_input[37088:37095] = '{32'hc276e6a1, 32'hc25d1502, 32'hc1f1b8c9, 32'hc09fc2d6, 32'h42990015, 32'hc074e0e4, 32'h41e90a29, 32'h41280366};
test_label[4636] = '{32'hc276e6a1};
test_output[4636] = '{32'h430a39b3};
/*############ DEBUG ############
test_input[37088:37095] = '{-61.7252233281, -55.2705166764, -30.2152275287, -4.99253369858, 76.5001629011, -3.82622631746, 29.1299616619, 10.5008299939};
test_label[4636] = '{-61.7252233281};
test_output[4636] = '{138.225386229};
############ END DEBUG ############*/
test_input[37096:37103] = '{32'h4214767f, 32'h428c9f03, 32'h41f61741, 32'hc09aef40, 32'hc2c550e4, 32'hc1356835, 32'hc1ccdd19, 32'h42898ab0};
test_label[4637] = '{32'h41f61741};
test_output[4637] = '{32'h421ef959};
/*############ DEBUG ############
test_input[37096:37103] = '{37.1157174882, 70.3105688126, 30.7613552988, -4.84170513847, -98.6579892249, -11.3379414469, -25.6079583868, 68.7708762046};
test_label[4637] = '{30.7613552988};
test_output[4637] = '{39.7435023516};
############ END DEBUG ############*/
test_input[37104:37111] = '{32'h42bd58a5, 32'h42a10fed, 32'h42aad2ce, 32'hc269fe82, 32'hc183fa30, 32'h42a9325e, 32'h42668cbf, 32'h423d7b2d};
test_label[4638] = '{32'h42aad2ce};
test_output[4638] = '{32'h41142f49};
/*############ DEBUG ############
test_input[37104:37111] = '{94.6731312727, 80.5311037434, 85.4117250117, -58.4985428559, -16.4971623796, 84.5983718735, 57.6374463588, 47.3702870487};
test_label[4638] = '{85.4117250117};
test_output[4638] = '{9.26154412414};
############ END DEBUG ############*/
test_input[37112:37119] = '{32'h42639bd1, 32'hc20a1770, 32'hc29358a2, 32'h41b99c1e, 32'hc29e18a8, 32'hc265f783, 32'h418fe635, 32'h41f4208e};
test_label[4639] = '{32'h41f4208e};
test_output[4639] = '{32'h41d31713};
/*############ DEBUG ############
test_input[37112:37119] = '{56.9021632339, -34.5228888527, -73.6731137968, 23.201229149, -79.0481567182, -57.4917113589, 17.9874061697, 30.5158962282};
test_label[4639] = '{30.5158962282};
test_output[4639] = '{26.3862670057};
############ END DEBUG ############*/
test_input[37120:37127] = '{32'h42bdcf80, 32'hc09de23c, 32'hc29d0d33, 32'hc2af39d8, 32'h4200d360, 32'hc174ef3f, 32'hc2427fc2, 32'hc281b2e2};
test_label[4640] = '{32'hc09de23c};
test_output[4640] = '{32'h42c7ada4};
/*############ DEBUG ############
test_input[37120:37127] = '{94.9052729982, -4.93386638642, -78.5257777417, -87.6129782994, 32.2064226163, -15.3084099056, -48.624764525, -64.8493837096};
test_label[4640] = '{-4.93386638642};
test_output[4640] = '{99.8391393846};
############ END DEBUG ############*/
test_input[37128:37135] = '{32'hc29a65e3, 32'h42675d27, 32'hc26af7cd, 32'hc26eba1e, 32'h423bd946, 32'h4299e6b1, 32'hc2a792b3, 32'h41ec6a8e};
test_label[4641] = '{32'hc2a792b3};
test_output[4641] = '{32'h4320bcb2};
/*############ DEBUG ############
test_input[37128:37135] = '{-77.1990001432, 57.8409689761, -58.7419914251, -59.6817548841, 46.9621802033, 76.9505707016, -83.7865189622, 29.5520283304};
test_label[4641] = '{-83.7865189622};
test_output[4641] = '{160.737089669};
############ END DEBUG ############*/
test_input[37136:37143] = '{32'h42849ba7, 32'h428545d9, 32'h429470d5, 32'hc28a71ba, 32'hc2195912, 32'h42852946, 32'h422a7461, 32'h4108887b};
test_label[4642] = '{32'h422a7461};
test_output[4642] = '{32'h41fcdd57};
/*############ DEBUG ############
test_input[37136:37143] = '{66.3040049532, 66.6364211713, 74.2203740896, -69.222125824, -38.3369840505, 66.580608697, 42.6136512637, 8.5333205357};
test_label[4642] = '{42.6136512637};
test_output[4642] = '{31.6080761222};
############ END DEBUG ############*/
test_input[37144:37151] = '{32'hc19eae9a, 32'h4289ad57, 32'h423601e2, 32'h418bae5b, 32'h42358076, 32'hc280839b, 32'hc2b6caec, 32'h42c68887};
test_label[4643] = '{32'h4289ad57};
test_output[4643] = '{32'h41f36cc1};
/*############ DEBUG ############
test_input[37144:37151] = '{-19.8352537592, 68.8385553505, 45.5018383404, 17.4601349722, 45.3754488468, -64.2570455186, -91.3963346057, 99.2666576179};
test_label[4643] = '{68.8385553505};
test_output[4643] = '{30.4281022675};
############ END DEBUG ############*/
test_input[37152:37159] = '{32'hc192eb0e, 32'h42876c50, 32'h42224126, 32'h4120f8b7, 32'hc252a604, 32'hc28ff8a9, 32'h41c7d3f3, 32'h4150e5bb};
test_label[4644] = '{32'h41c7d3f3};
test_output[4644] = '{32'h422aeea7};
/*############ DEBUG ############
test_input[37152:37159] = '{-18.3647719379, 67.7115476149, 40.5636210724, 10.0607212135, -52.6621231501, -71.9856629352, 24.978490285, 13.0560862522};
test_label[4644] = '{24.978490285};
test_output[4644] = '{42.7330573298};
############ END DEBUG ############*/
test_input[37160:37167] = '{32'hc157e607, 32'h41c416f9, 32'hc20dfebe, 32'hc2c6335c, 32'h4293be1a, 32'h423cdb06, 32'hc2b008a7, 32'hbf1d00e7};
test_label[4645] = '{32'hc20dfebe};
test_output[4645] = '{32'h42dabd79};
/*############ DEBUG ############
test_input[37160:37167] = '{-13.4936589541, 24.5112163098, -35.4987724872, -99.1003122404, 73.871292325, 47.2138899369, -88.0169006012, -0.613295001954};
test_label[4645] = '{-35.4987724872};
test_output[4645] = '{109.370064812};
############ END DEBUG ############*/
test_input[37168:37175] = '{32'h4296df98, 32'h429a725b, 32'h40de8ef7, 32'h426c05d9, 32'h416943f9, 32'h425ad850, 32'h40da8c10, 32'h40aeebb8};
test_label[4646] = '{32'h426c05d9};
test_output[4646] = '{32'h4192faec};
/*############ DEBUG ############
test_input[37168:37175] = '{75.4367030543, 77.2233468039, 6.95495193779, 59.0057097358, 14.5790944486, 54.7112435614, 6.82959758784, 5.4662741501};
test_label[4646] = '{59.0057097358};
test_output[4646] = '{18.3725201798};
############ END DEBUG ############*/
test_input[37176:37183] = '{32'h412d9a5d, 32'hc22a5a5f, 32'h42864fd8, 32'hc1ce9230, 32'hc18167df, 32'h425f371c, 32'h420da112, 32'h41dd9f82};
test_label[4647] = '{32'h41dd9f82};
test_output[4647] = '{32'h421dcff2};
/*############ DEBUG ############
test_input[37176:37183] = '{10.8501860862, -42.5882541972, 67.1559451696, -25.8213810792, -16.1757184517, 55.8038170829, 35.4072970505, 27.7028854102};
test_label[4647] = '{27.7028854102};
test_output[4647] = '{39.4530715039};
############ END DEBUG ############*/
test_input[37184:37191] = '{32'h41dd0d18, 32'hc290d9e4, 32'h4014e9b3, 32'h42c2e3b3, 32'h42a253ca, 32'h42bf7ca4, 32'hc29f082f, 32'hc2b0ad58};
test_label[4648] = '{32'hc290d9e4};
test_output[4648] = '{32'h432a09b2};
/*############ DEBUG ############
test_input[37184:37191] = '{27.6313936931, -72.4255673866, 2.32676398621, 97.4447226437, 81.1636518478, 95.7434358532, -79.5159819059, -88.3385603772};
test_label[4648] = '{-72.4255673866};
test_output[4648] = '{170.037877475};
############ END DEBUG ############*/
test_input[37192:37199] = '{32'h40cc218c, 32'h41a9e06e, 32'h424ff3bb, 32'hc0d63840, 32'hc27a7778, 32'hc0925ca0, 32'hc2b5028a, 32'h4268acda};
test_label[4649] = '{32'hc2b5028a};
test_output[4649] = '{32'h4314ad03};
/*############ DEBUG ############
test_input[37192:37199] = '{6.37909489484, 21.2345846756, 51.9880184047, -6.69436662122, -62.6166700023, -4.57380698457, -90.5049627635, 58.1688003522};
test_label[4649] = '{-90.5049627635};
test_output[4649] = '{148.675829788};
############ END DEBUG ############*/
test_input[37200:37207] = '{32'hc2737ef0, 32'hc096f6ab, 32'h4266699d, 32'hc2a16ee6, 32'h42359c27, 32'h422d256b, 32'hc297c439, 32'h42ba0415};
test_label[4650] = '{32'h42359c27};
test_output[4650] = '{32'h423e6c02};
/*############ DEBUG ############
test_input[37200:37207] = '{-60.8739622037, -4.7176109171, 57.6031380564, -80.7165965361, 45.4024929318, 43.2865422188, -75.8832474646, 93.0079697042};
test_label[4650] = '{45.4024929318};
test_output[4650] = '{47.6054767724};
############ END DEBUG ############*/
test_input[37208:37215] = '{32'hc2729751, 32'h429f151b, 32'h42aec3bc, 32'h41ff15cf, 32'hc2bdfa48, 32'h429c60d6, 32'hc2014e86, 32'h424c2a68};
test_label[4651] = '{32'hc2014e86};
test_output[4651] = '{32'h42ef6b40};
/*############ DEBUG ############
test_input[37208:37215] = '{-60.6477711193, 79.5412225174, 87.382291527, 31.8856479717, -94.9888315802, 78.1891322954, -32.326683782, 51.0414115693};
test_label[4651] = '{-32.326683782};
test_output[4651] = '{119.709470168};
############ END DEBUG ############*/
test_input[37216:37223] = '{32'hc1804c2d, 32'h42693edc, 32'h4288c1ac, 32'hc1eded44, 32'h40b32bb9, 32'h420a5526, 32'hc1c68033, 32'hc252ddcb};
test_label[4652] = '{32'h40b32bb9};
test_output[4652] = '{32'h427b1deb};
/*############ DEBUG ############
test_input[37216:37223] = '{-16.0371953716, 58.3113849471, 68.3782630141, -29.7408528776, 5.59908725919, 34.5831528462, -24.8125972982, -52.7165945626};
test_label[4652] = '{5.59908725919};
test_output[4652] = '{62.779218217};
############ END DEBUG ############*/
test_input[37224:37231] = '{32'hc14b7a25, 32'h42079ba9, 32'hc1eb31a0, 32'hc2a05b52, 32'h424d404d, 32'h40a46b38, 32'hc22ad702, 32'h42a82286};
test_label[4653] = '{32'h424d404d};
test_output[4653] = '{32'h420304bf};
/*############ DEBUG ############
test_input[37224:37231] = '{-12.7173206872, 33.9020117347, -29.3992318093, -80.1783613808, 51.3127952543, 5.13808805554, -42.7099701521, 84.0674308227};
test_label[4653] = '{51.3127952543};
test_output[4653] = '{32.7546355683};
############ END DEBUG ############*/
test_input[37232:37239] = '{32'hc291185e, 32'h40b91fed, 32'h404a5b18, 32'h41f803de, 32'hc226345c, 32'h3f4751ed, 32'h42ab8eb5, 32'h428a1b8a};
test_label[4654] = '{32'h428a1b8a};
test_output[4654] = '{32'h4185ccab};
/*############ DEBUG ############
test_input[37232:37239] = '{-72.5475947429, 5.78514737893, 3.16180991069, 31.0018889896, -41.5511319163, 0.778593862632, 85.778724534, 69.0537885197};
test_label[4654] = '{69.0537885197};
test_output[4654] = '{16.7249360689};
############ END DEBUG ############*/
test_input[37240:37247] = '{32'h41f92937, 32'hc151e1b8, 32'hc14bb72a, 32'hc230d4b3, 32'hc1f60247, 32'hc21c14a3, 32'hc23419ec, 32'h423170b5};
test_label[4655] = '{32'hc14bb72a};
test_output[4655] = '{32'h42645e80};
/*############ DEBUG ############
test_input[37240:37247] = '{31.1451248398, -13.1176070737, -12.7322179794, -44.2077158301, -30.7511116268, -39.0201526031, -45.0253133898, 44.3600647827};
test_label[4655] = '{-12.7322179794};
test_output[4655] = '{57.0922845853};
############ END DEBUG ############*/
test_input[37248:37255] = '{32'h427d6581, 32'h41ab62b0, 32'h42bfa65d, 32'h42af67dd, 32'h4195ee81, 32'h4271666d, 32'hc2b5fcb5, 32'hc266b4b7};
test_label[4656] = '{32'h4195ee81};
test_output[4656] = '{32'h429a2ae3};
/*############ DEBUG ############
test_input[37248:37255] = '{63.3491256406, 21.4231879363, 95.8249264094, 87.7028563291, 18.7414571425, 60.3500243156, -90.9935647234, -57.6764795363};
test_label[4656] = '{18.7414571425};
test_output[4656] = '{77.0837661362};
############ END DEBUG ############*/
test_input[37256:37263] = '{32'h428fcc0c, 32'h408c1f24, 32'h428efecf, 32'hc28f089c, 32'hc205d001, 32'h4108cfa8, 32'h42adab48, 32'hc2782a51};
test_label[4657] = '{32'hc2782a51};
test_output[4657] = '{32'h4314e038};
/*############ DEBUG ############
test_input[37256:37263] = '{71.8985276826, 4.37880150273, 71.4976714089, -71.5168182363, -33.4531284321, 8.55069730161, 86.8345314597, -62.0413256802};
test_label[4657] = '{-62.0413256802};
test_output[4657] = '{148.875857684};
############ END DEBUG ############*/
test_input[37264:37271] = '{32'h411a6074, 32'h3e8cd0ef, 32'h42abdd4a, 32'h4228df2a, 32'h4209581d, 32'h429f42f0, 32'h42be7936, 32'h40b00637};
test_label[4658] = '{32'h4209581d};
test_output[4658] = '{32'h42739a67};
/*############ DEBUG ############
test_input[37264:37271] = '{9.64854781149, 0.275031549639, 85.9322047659, 42.217934134, 34.3360476434, 79.6307377169, 95.2367401831, 5.5007585117};
test_label[4658] = '{34.3360476434};
test_output[4658] = '{60.9007837129};
############ END DEBUG ############*/
test_input[37272:37279] = '{32'hc2182e6f, 32'hc2377d07, 32'h41597488, 32'h423d023b, 32'h408b4c93, 32'h3f8bec15, 32'hc20f91b4, 32'hc076685c};
test_label[4659] = '{32'h41597488};
test_output[4659] = '{32'h4206a519};
/*############ DEBUG ############
test_input[37272:37279] = '{-38.0453446099, -45.8720971565, 13.590949874, 47.2521777964, 4.35309738168, 1.09314218748, -35.8922873283, -3.85011970937};
test_label[4659] = '{13.590949874};
test_output[4659] = '{33.6612279224};
############ END DEBUG ############*/
test_input[37280:37287] = '{32'h420d6b74, 32'h42bdbb02, 32'h401c3501, 32'h42a24ed5, 32'h419fec0e, 32'h421a1ea0, 32'h420542fd, 32'h411ea30a};
test_label[4660] = '{32'h42a24ed5};
test_output[4660] = '{32'h415b616d};
/*############ DEBUG ############
test_input[37280:37287] = '{35.3549336764, 94.8652505681, 2.440734996, 81.1539660364, 19.990261302, 38.5299071178, 33.3154176092, 9.91480482496};
test_label[4660] = '{81.1539660364};
test_output[4660] = '{13.7112856416};
############ END DEBUG ############*/
test_input[37288:37295] = '{32'h4246223f, 32'h4243eb85, 32'hc15327b2, 32'h428e88ce, 32'hc1b8ea11, 32'h418d5743, 32'hc23e7b4e, 32'hc2a2b858};
test_label[4661] = '{32'h418d5743};
test_output[4661] = '{32'h425665fa};
/*############ DEBUG ############
test_input[37288:37295] = '{49.5334425806, 48.980000366, -13.197191642, 71.267194732, -23.1142904092, 17.6676089464, -47.6204162776, -81.3600472764};
test_label[4661] = '{17.6676089464};
test_output[4661] = '{53.5995857861};
############ END DEBUG ############*/
test_input[37296:37303] = '{32'h4269a5d7, 32'hc2a4a8a3, 32'h414027c1, 32'h41a723bb, 32'hc133eaa1, 32'h42556fce, 32'h3f8387de, 32'hc09e64b7};
test_label[4662] = '{32'h414027c1};
test_output[4662] = '{32'h4239a26d};
/*############ DEBUG ############
test_input[37296:37303] = '{58.4119541612, -82.3293653155, 12.0097059954, 20.8924459854, -11.2447829051, 53.3591848764, 1.02758381461, -4.94979411108};
test_label[4662] = '{12.0097059954};
test_output[4662] = '{46.4086194348};
############ END DEBUG ############*/
test_input[37304:37311] = '{32'h429af787, 32'h4258f463, 32'hc2a6f97c, 32'hc284c3e2, 32'h402e2169, 32'h422aa42c, 32'h41c5f6bb, 32'h4242300d};
test_label[4663] = '{32'h41c5f6bb};
test_output[4663] = '{32'h4252f3b1};
/*############ DEBUG ############
test_input[37304:37311] = '{77.4834545122, 54.238658472, -83.4872739595, -66.382581507, 2.7207891122, 42.6603257062, 24.7454740998, 48.5469254528};
test_label[4663] = '{24.7454740998};
test_output[4663] = '{52.7379804125};
############ END DEBUG ############*/
test_input[37312:37319] = '{32'h4228122f, 32'h4212b12c, 32'h4272f3ec, 32'h415e345c, 32'h427002ab, 32'h4100a8b3, 32'hc205b17b, 32'hc2850a72};
test_label[4664] = '{32'h427002ab};
test_output[4664] = '{32'h3f904542};
/*############ DEBUG ############
test_input[37312:37319] = '{42.0177569143, 36.6730184777, 60.7382067165, 13.8877829784, 60.0026064674, 8.04118671013, -33.4233192777, -66.5204001007};
test_label[4664] = '{60.0026064674};
test_output[4664] = '{1.12711363636};
############ END DEBUG ############*/
test_input[37320:37327] = '{32'h41603aa9, 32'hc2baeca5, 32'hc22b08a8, 32'h4296f2f8, 32'hc08ce728, 32'h41a018b0, 32'h413cd6e2, 32'hc2b1bfe2};
test_label[4665] = '{32'hc2b1bfe2};
test_output[4665] = '{32'h4324596d};
/*############ DEBUG ############
test_input[37320:37327] = '{14.0143210057, -93.4621940362, -42.7584547063, 75.4745455034, -4.40321713722, 20.0120546139, 11.802461296, -88.8747724252};
test_label[4665] = '{-88.8747724252};
test_output[4665] = '{164.349317929};
############ END DEBUG ############*/
test_input[37328:37335] = '{32'h423f253d, 32'h41cd0667, 32'h42008cd7, 32'h415d1380, 32'hc28fe776, 32'hc2c636fa, 32'hc2b36e25, 32'hc2383396};
test_label[4666] = '{32'h42008cd7};
test_output[4666] = '{32'h417a6198};
/*############ DEBUG ############
test_input[37328:37335] = '{47.7863663114, 25.6281257928, 32.1375397008, 13.8172610886, -71.9520707113, -99.1073789297, -89.7151261658, -46.0503782042};
test_label[4666] = '{32.1375397008};
test_output[4666] = '{15.6488267707};
############ END DEBUG ############*/
test_input[37336:37343] = '{32'h4222c534, 32'hc22bc8ad, 32'hc187d9db, 32'hc13ddf03, 32'h42b8ae72, 32'h41a261ba, 32'h42968d6e, 32'h4045b9fb};
test_label[4667] = '{32'h4222c534};
test_output[4667] = '{32'h424e97af};
/*############ DEBUG ############
test_input[37336:37343] = '{40.6925817021, -42.9459737679, -16.9813742562, -11.8669461815, 92.3407099522, 20.2977171205, 75.2762326194, 3.08947645258};
test_label[4667] = '{40.6925817021};
test_output[4667] = '{51.6481282889};
############ END DEBUG ############*/
test_input[37344:37351] = '{32'hc15b678c, 32'hc271000c, 32'hc2204e14, 32'h4280ea71, 32'hc20ea697, 32'hc2aea3fa, 32'h419080a4, 32'h429facd6};
test_label[4668] = '{32'hc20ea697};
test_output[4668] = '{32'h42e70022};
/*############ DEBUG ############
test_input[37344:37351] = '{-13.7127798194, -60.2500448455, -40.0762470626, 64.4578915198, -35.6626867274, -87.3202673583, 18.0628126291, 79.8375725968};
test_label[4668] = '{-35.6626867274};
test_output[4668] = '{115.500259533};
############ END DEBUG ############*/
test_input[37352:37359] = '{32'h42593ca5, 32'hc231d7a3, 32'h42a0aa9f, 32'hc2185971, 32'h42a9320b, 32'h42b7222d, 32'hc12fe27d, 32'h423d5653};
test_label[4669] = '{32'h423d5653};
test_output[4669] = '{32'h4230ef01};
/*############ DEBUG ############
test_input[37352:37359] = '{54.3092224561, -44.460584373, 80.3332465045, -38.0873436995, 84.5977406088, 91.5667471693, -10.9927952089, 47.3342993621};
test_label[4669] = '{47.3342993621};
test_output[4669] = '{44.2334011631};
############ END DEBUG ############*/
test_input[37360:37367] = '{32'hc197b792, 32'hc21de4af, 32'hc1ae73ab, 32'hc29c2502, 32'hc27d0e1a, 32'hc2817b12, 32'hc1441dcf, 32'hc2691165};
test_label[4670] = '{32'hc2817b12};
test_output[4670] = '{32'h4251f003};
/*############ DEBUG ############
test_input[37360:37367] = '{-18.9646346097, -39.4733241605, -21.8064777696, -78.0722842994, -63.263772483, -64.7403701403, -12.257277743, -58.266985836};
test_label[4670] = '{-64.7403701403};
test_output[4670] = '{52.4843847096};
############ END DEBUG ############*/
test_input[37368:37375] = '{32'h41f06b65, 32'h428fe19e, 32'h3f8ac88b, 32'hc2b4b1c9, 32'h428efb3f, 32'hc24114ad, 32'h419880d4, 32'h4297c126};
test_label[4671] = '{32'hc24114ad};
test_output[4671] = '{32'h42f85b98};
/*############ DEBUG ############
test_input[37368:37375] = '{30.0524391409, 71.9406618315, 1.08424505813, -90.3472395307, 71.4907132537, -48.2701917557, 19.0629045632, 75.8772438688};
test_label[4671] = '{-48.2701917557};
test_output[4671] = '{124.178894202};
############ END DEBUG ############*/
test_input[37376:37383] = '{32'hc08a535e, 32'hbfd4a8de, 32'hc2aaa8e8, 32'hc2b08e4a, 32'hc21ea780, 32'h41346152, 32'hc2924683, 32'hc2916506};
test_label[4672] = '{32'hbfd4a8de};
test_output[4672] = '{32'h414ef670};
/*############ DEBUG ############
test_input[37376:37383] = '{-4.32267655206, -1.66140347451, -85.3298983216, -88.2779071031, -39.663574395, 11.273759412, -73.1377188212, -72.6973102914};
test_label[4672] = '{-1.66140347451};
test_output[4672] = '{12.9351654668};
############ END DEBUG ############*/
test_input[37384:37391] = '{32'hc23e2765, 32'hc26613be, 32'h42841d6b, 32'hc1fa89cd, 32'hc2341195, 32'h41da11eb, 32'h4221a1c4, 32'hc20d49bc};
test_label[4673] = '{32'hc20d49bc};
test_output[4673] = '{32'h42cac249};
/*############ DEBUG ############
test_input[37384:37391] = '{-47.5384727862, -57.5192809553, 66.0574600038, -31.3172849572, -45.0171681894, 27.2587498637, 40.4079744944, -35.3220054549};
test_label[4673] = '{-35.3220054549};
test_output[4673] = '{101.379465459};
############ END DEBUG ############*/
test_input[37392:37399] = '{32'hc234cb3c, 32'hc14b6f5c, 32'h423b5780, 32'h429d229c, 32'h420678f6, 32'hc21a6b20, 32'hc2374f42, 32'h421f109b};
test_label[4674] = '{32'h423b5780};
test_output[4674] = '{32'h41fddb71};
/*############ DEBUG ############
test_input[37392:37399] = '{-45.198469628, -12.7146876786, 46.8354503978, 78.5675993714, 33.6181263583, -38.6046133987, -45.8274014144, 39.7662145946};
test_label[4674] = '{46.8354503978};
test_output[4674] = '{31.7321489736};
############ END DEBUG ############*/
test_input[37400:37407] = '{32'h42c56984, 32'h42a81f46, 32'h4234c3eb, 32'h42999e24, 32'h4252c541, 32'h4261e961, 32'hc285cb5e, 32'hc27a8665};
test_label[4675] = '{32'h4261e961};
test_output[4675] = '{32'h4228e9a7};
/*############ DEBUG ############
test_input[37400:37407] = '{98.7060850836, 84.0610778947, 45.1913279359, 76.8088661883, 52.6926297302, 56.4779093035, -66.8972051729, -62.6312431644};
test_label[4675] = '{56.4779093035};
test_output[4675] = '{42.2281762167};
############ END DEBUG ############*/
test_input[37408:37415] = '{32'hc2a196bd, 32'h41a508ad, 32'hc14b5e77, 32'hc24b2e3e, 32'hc2955d64, 32'hc1b842e8, 32'h42bcb6f5, 32'h41cb5feb};
test_label[4676] = '{32'h41cb5feb};
test_output[4676] = '{32'h4289defa};
/*############ DEBUG ############
test_input[37408:37415] = '{-80.794411832, 20.6292361248, -12.7105630381, -50.7951567347, -74.6824028466, -23.0326691586, 94.3573398762, 25.4218352146};
test_label[4676] = '{25.4218352146};
test_output[4676] = '{68.9355046615};
############ END DEBUG ############*/
test_input[37416:37423] = '{32'hc1814806, 32'hc2abf39b, 32'h42ad1eae, 32'h41b5b50c, 32'hc28657f5, 32'h41bf9e14, 32'hc2536880, 32'h424ec500};
test_label[4677] = '{32'hc28657f5};
test_output[4677] = '{32'h4319bb51};
/*############ DEBUG ############
test_input[37416:37423] = '{-16.1601681089, -85.9757882002, 86.5599186506, 22.7134018805, -67.1717909806, 23.9521868603, -52.8520506358, 51.6923812107};
test_label[4677] = '{-67.1717909806};
test_output[4677] = '{153.731709631};
############ END DEBUG ############*/
test_input[37424:37431] = '{32'h41abc334, 32'h42647c68, 32'hc18577a8, 32'h4282d039, 32'hc1ff1c5d, 32'hc285c915, 32'h414fe45c, 32'h42bb6a82};
test_label[4678] = '{32'h414fe45c};
test_output[4678] = '{32'h42a16df7};
/*############ DEBUG ############
test_input[37424:37431] = '{21.4703136873, 57.1214904373, -16.6834254323, 65.4066864095, -31.8888491668, -66.8927351236, 12.993251681, 93.7080247307};
test_label[4678] = '{12.993251681};
test_output[4678] = '{80.7147730497};
############ END DEBUG ############*/
test_input[37432:37439] = '{32'hc2772ca1, 32'h4183084e, 32'h41e624d4, 32'hc2a93cc1, 32'h424c58ae, 32'hc10dea43, 32'hc15012fe, 32'h42559f6e};
test_label[4679] = '{32'h41e624d4};
test_output[4679] = '{32'h41c5da2d};
/*############ DEBUG ############
test_input[37432:37439] = '{-61.7935840587, 16.3790549201, 28.7679833428, -84.6186628759, 51.086599399, -8.86969323535, -13.0046371082, 53.4056929511};
test_label[4679] = '{28.7679833428};
test_output[4679] = '{24.73153023};
############ END DEBUG ############*/
test_input[37440:37447] = '{32'hc294322b, 32'hc1ad47ec, 32'h41c947d5, 32'h41d16d90, 32'hc2ab7c5e, 32'h424de51c, 32'hc2c3b4e4, 32'h4261b7b2};
test_label[4680] = '{32'h4261b7b2};
test_output[4680] = '{32'h3be5fe33};
/*############ DEBUG ############
test_input[37440:37447] = '{-74.0979847346, -21.6601176731, 25.1600738235, 26.1784970837, -85.7429074412, 51.4737414592, -97.8533039588, 56.4293890012};
test_label[4680] = '{56.4293890012};
test_output[4680] = '{0.00701882812489};
############ END DEBUG ############*/
test_input[37448:37455] = '{32'h4298266c, 32'hc2c694f5, 32'h3f878259, 32'hc189ebb9, 32'hc0875a42, 32'h429e5504, 32'hc2b82168, 32'h4236935d};
test_label[4681] = '{32'hc0875a42};
test_output[4681] = '{32'h42a6e16b};
/*############ DEBUG ############
test_input[37448:37455] = '{76.0750415219, -99.2909331178, 1.0586654342, -17.2400992205, -4.22976797121, 79.1660499225, -92.0652464477, 45.6439105628};
test_label[4681] = '{-4.22976797121};
test_output[4681] = '{83.4402711369};
############ END DEBUG ############*/
test_input[37456:37463] = '{32'h424037a3, 32'hc1a09227, 32'h41f4d973, 32'hc2b75d84, 32'h41c7927d, 32'hbfa5620a, 32'h42b53233, 32'hc23c078a};
test_label[4682] = '{32'hc23c078a};
test_output[4682] = '{32'h43099afc};
/*############ DEBUG ############
test_input[37456:37463] = '{48.0543346396, -20.0713637591, 30.6061759376, -91.6826465824, 24.9465266903, -1.29205442217, 90.5980476402, -47.0073640253};
test_label[4682] = '{-47.0073640253};
test_output[4682] = '{137.605411665};
############ END DEBUG ############*/
test_input[37464:37471] = '{32'h422075c0, 32'h41a00d0b, 32'hc19b27d0, 32'h42b47a0a, 32'h428b6fbc, 32'hc1d48800, 32'h420bdd50, 32'hc2652d24};
test_label[4683] = '{32'h428b6fbc};
test_output[4683] = '{32'h41a42935};
/*############ DEBUG ############
test_input[37464:37471] = '{40.1149901553, 20.0063677416, -19.3944397411, 90.2383552656, 69.718234526, -26.5664064857, 34.9661267261, -57.2940814775};
test_label[4683] = '{69.718234526};
test_output[4683] = '{20.5201207409};
############ END DEBUG ############*/
test_input[37472:37479] = '{32'hc2967f26, 32'hc211ff35, 32'h426d9c5d, 32'hc2c6bd63, 32'hc225a554, 32'hc2b7d5eb, 32'h420eae50, 32'hc2b02699};
test_label[4684] = '{32'hc2b02699};
test_output[4684] = '{32'h43137a64};
/*############ DEBUG ############
test_input[37472:37479] = '{-75.2483405737, -36.4992249358, 59.40269763, -99.3698967023, -41.4114546601, -91.9178100519, 35.6702289075, -88.0753851496};
test_label[4684] = '{-88.0753851496};
test_output[4684] = '{147.47808278};
############ END DEBUG ############*/
test_input[37480:37487] = '{32'h4126ab2f, 32'hc25ac2aa, 32'h40c2feff, 32'h4212889c, 32'hc2996db1, 32'hc2a6c1f1, 32'hc210f1c3, 32'hc289c18e};
test_label[4685] = '{32'hc2a6c1f1};
test_output[4685] = '{32'h42f0063f};
/*############ DEBUG ############
test_input[37480:37487] = '{10.4167928999, -54.6901007759, 6.09362757677, 36.6334082419, -76.7142382604, -83.3787904871, -36.2360957385, -68.8780364268};
test_label[4685] = '{-83.3787904871};
test_output[4685] = '{120.012198729};
############ END DEBUG ############*/
test_input[37488:37495] = '{32'h4187d7d1, 32'hc2b1dc6a, 32'h42b7c96c, 32'hc1a19ff0, 32'hc29d7354, 32'hc2ad88bf, 32'hc1a489d3, 32'h42adbc7e};
test_label[4686] = '{32'hc29d7354};
test_output[4686] = '{32'h432aa00d};
/*############ DEBUG ############
test_input[37488:37495] = '{16.980379877, -88.93049505, 91.8934031676, -20.2030936945, -78.725249737, -86.767080205, -20.5672964399, 86.8681504871};
test_label[4686] = '{-78.725249737};
test_output[4686] = '{170.625201343};
############ END DEBUG ############*/
test_input[37496:37503] = '{32'h428e2f8a, 32'hc294e4e9, 32'h4293409a, 32'hc2034290, 32'h42b35897, 32'hc2a8ad78, 32'hc1fd1a85, 32'h413c823c};
test_label[4687] = '{32'hc2a8ad78};
test_output[4687] = '{32'h432e0308};
/*############ DEBUG ############
test_input[37496:37503] = '{71.0928496929, -74.4470891197, 73.6261747974, -32.8150032902, 89.6730243393, -84.3388088883, -31.6379487359, 11.7817952901};
test_label[4687] = '{-84.3388088883};
test_output[4687] = '{174.011833344};
############ END DEBUG ############*/
test_input[37504:37511] = '{32'hc28aac28, 32'h4261db2e, 32'hc2c5a9d0, 32'hc2b28ac9, 32'hc1955ebd, 32'h42c1ffc9, 32'h42c7d5fd, 32'hc29527bb};
test_label[4688] = '{32'hc29527bb};
test_output[4688] = '{32'h432e8c54};
/*############ DEBUG ############
test_input[37504:37511] = '{-69.3362388997, 56.4640442093, -98.8316680923, -89.2710627003, -18.6712593338, 96.9995841543, 99.9179457913, -74.5776018424};
test_label[4688] = '{-74.5776018424};
test_output[4688] = '{174.548161073};
############ END DEBUG ############*/
test_input[37512:37519] = '{32'h41f685a8, 32'hc1e99a92, 32'hc2766d2f, 32'hc23109b2, 32'hc233f0e4, 32'h416298a6, 32'hc2227b83, 32'h419a7cf2};
test_label[4689] = '{32'hc233f0e4};
test_output[4689] = '{32'h429799dd};
/*############ DEBUG ############
test_input[37512:37519] = '{30.8152612349, -29.2004730395, -61.606625778, -44.259466412, -44.9852464734, 14.162267614, -40.6206167136, 19.3110090949};
test_label[4689] = '{-44.9852464734};
test_output[4689] = '{75.8005178539};
############ END DEBUG ############*/
test_input[37520:37527] = '{32'hc2af9574, 32'h421458d8, 32'h41af40b0, 32'hc2401dd0, 32'h4290f99b, 32'h41bec147, 32'hc29197a6, 32'h4235133d};
test_label[4690] = '{32'h41af40b0};
test_output[4690] = '{32'h424a52de};
/*############ DEBUG ############
test_input[37520:37527] = '{-87.7919026158, 37.0867612757, 21.906585569, -48.0291120337, 72.4875093559, 23.8443739072, -72.7961901622, 45.2687881335};
test_label[4690] = '{21.906585569};
test_output[4690] = '{50.5809237869};
############ END DEBUG ############*/
test_input[37528:37535] = '{32'h421758b6, 32'hc28e20a8, 32'hc258897d, 32'h41f123ee, 32'h421a745b, 32'h425223ff, 32'hc2876518, 32'h41a843ff};
test_label[4691] = '{32'hc28e20a8};
test_output[4691] = '{32'h42f732a8};
/*############ DEBUG ############
test_input[37528:37535] = '{37.8366299675, -71.0637817225, -54.1342641775, 30.1425437351, 38.6136288705, 52.5351513584, -67.6974510736, 21.0332021007};
test_label[4691] = '{-71.0637817225};
test_output[4691] = '{123.598934394};
############ END DEBUG ############*/
test_input[37536:37543] = '{32'h420c4598, 32'hc2a53e32, 32'h41c63994, 32'hc282c5e6, 32'h40dc0d42, 32'h42b81376, 32'hc17a8678, 32'hc285499b};
test_label[4692] = '{32'hc285499b};
test_output[4692] = '{32'h431eae88};
/*############ DEBUG ############
test_input[37536:37543] = '{35.067962314, -82.6214738436, 24.7781145427, -65.3865232985, 6.87661854792, 92.0380060408, -15.6578296848, -66.6437597246};
test_label[4692] = '{-66.6437597246};
test_output[4692] = '{158.681765765};
############ END DEBUG ############*/
test_input[37544:37551] = '{32'hc04032de, 32'h4227dff2, 32'hc2953caa, 32'h41f4ff36, 32'hc21c1376, 32'h42869efb, 32'hc1a77d7d, 32'hc1e19962};
test_label[4693] = '{32'hc1e19962};
test_output[4693] = '{32'h42bf0553};
/*############ DEBUG ############
test_input[37544:37551] = '{-3.00310465645, 41.9686961942, -74.6184848434, 30.62461478, -39.0190066294, 67.3105057285, -20.9362737996, -28.1998930476};
test_label[4693] = '{-28.1998930476};
test_output[4693] = '{95.5103987762};
############ END DEBUG ############*/
test_input[37552:37559] = '{32'hc1d49199, 32'h42a5f5ac, 32'h42211324, 32'hc0ce8d29, 32'hc236e149, 32'hc2261158, 32'hc2ba5f74, 32'hc173179b};
test_label[4694] = '{32'hc0ce8d29};
test_output[4694] = '{32'h42b2de7f};
/*############ DEBUG ############
test_input[37552:37559] = '{-26.5710931579, 82.9798300758, 40.2686919495, -6.45473135563, -45.720003561, -41.5169358847, -93.186428348, -15.193262833};
test_label[4694] = '{-6.45473135563};
test_output[4694] = '{89.4345614314};
############ END DEBUG ############*/
test_input[37560:37567] = '{32'hc28f483e, 32'h42132353, 32'hc105a8c7, 32'h3f9976c0, 32'h42876494, 32'hc29b756c, 32'hc11c9c02, 32'hc217614c};
test_label[4695] = '{32'hc105a8c7};
test_output[4695] = '{32'h429819ad};
/*############ DEBUG ############
test_input[37560:37567] = '{-71.6410965122, 36.7844961379, -8.35370525369, 1.19893642591, 67.696441753, -77.7293409929, -9.788087748, -37.8450172149};
test_label[4695] = '{-8.35370525369};
test_output[4695] = '{76.0501470067};
############ END DEBUG ############*/
test_input[37568:37575] = '{32'h42a4dc17, 32'h41b789a9, 32'h422ef3e7, 32'h426d3090, 32'hc2baeadc, 32'h42aa57a7, 32'h4134f2ae, 32'h41a9873d};
test_label[4696] = '{32'h422ef3e7};
test_output[4696] = '{32'h4225fb64};
/*############ DEBUG ############
test_input[37568:37575] = '{82.4298654945, 22.9422173184, 43.7381840948, 59.2974238724, -93.4587087228, 85.1711926043, 11.3092484428, 21.191035226};
test_label[4696] = '{43.7381840948};
test_output[4696] = '{41.4954993529};
############ END DEBUG ############*/
test_input[37576:37583] = '{32'h422d5f6f, 32'hc188f4b2, 32'h410c42d9, 32'hc0a129e6, 32'h41f62abe, 32'hc245a3ad, 32'h41b3956c, 32'hc25756d5};
test_label[4697] = '{32'h41f62abe};
test_output[4697] = '{32'h41492845};
/*############ DEBUG ############
test_input[37576:37583] = '{43.3431977507, -17.1194793826, 8.76632034131, -5.03636451718, 30.7708693565, -49.4098400734, 22.4479595044, -53.8347984404};
test_label[4697] = '{30.7708693565};
test_output[4697] = '{12.5723318617};
############ END DEBUG ############*/
test_input[37584:37591] = '{32'hc2327343, 32'hc20990a8, 32'h41e5f8c1, 32'hc24905ce, 32'h418e26d8, 32'hc20b9a91, 32'hc2b249b9, 32'h41a7071c};
test_label[4698] = '{32'h41e5f8c1};
test_output[4698] = '{32'h39d19ccf};
/*############ DEBUG ############
test_input[37584:37591] = '{-44.6125591558, -34.3912651036, 28.7464625959, -50.2556678484, 17.7689663097, -34.9009430995, -89.1439888182, 20.8784707216};
test_label[4698] = '{28.7464625959};
test_output[4698] = '{0.000399804185678};
############ END DEBUG ############*/
test_input[37592:37599] = '{32'h4295ff12, 32'h42b574bc, 32'hc250ac15, 32'h4141f14f, 32'h41d290e0, 32'hc2bebe08, 32'h42b9df7e, 32'h41257c5a};
test_label[4699] = '{32'hc250ac15};
test_output[4699] = '{32'h43113574};
/*############ DEBUG ############
test_input[37592:37599] = '{74.9981816989, 90.7279991966, -52.1680478327, 12.1214130986, 26.3207395028, -95.3711575657, 92.9365080994, 10.3428595112};
test_label[4699] = '{-52.1680478327};
test_output[4699] = '{145.208793743};
############ END DEBUG ############*/
test_input[37600:37607] = '{32'h41899b7c, 32'hc269fc79, 32'hc201fe84, 32'h42c56f08, 32'hc257047a, 32'hc2bc520d, 32'h41fafe76, 32'hc25aeeff};
test_label[4700] = '{32'hc269fc79};
test_output[4700] = '{32'h431d36a2};
/*############ DEBUG ############
test_input[37600:37607] = '{17.2009207728, -58.4965551597, -32.4985490354, 98.7168555725, -53.7543733777, -94.1602521764, 31.3742491356, -54.7333933288};
test_label[4700] = '{-58.4965551597};
test_output[4700] = '{157.213410732};
############ END DEBUG ############*/
test_input[37608:37615] = '{32'hc2aaaeb4, 32'hc23ad2b6, 32'hc295f853, 32'h4182cdde, 32'h4153e13d, 32'hc18a98ab, 32'hc1ee2163, 32'h3f07b83c};
test_label[4701] = '{32'hc18a98ab};
test_output[4701] = '{32'h4206e009};
/*############ DEBUG ############
test_input[37608:37615] = '{-85.3412198964, -46.7057724721, -74.9850100675, 16.3505207364, 13.2424895548, -17.3245453961, -29.7663012988, 0.530154950998};
test_label[4701] = '{-17.3245453961};
test_output[4701] = '{33.7187853542};
############ END DEBUG ############*/
test_input[37616:37623] = '{32'hc28d51dd, 32'h42bcb45c, 32'hc26816aa, 32'h42bb37aa, 32'hc28d95cc, 32'hc2af593a, 32'hc0505944, 32'h4184d2f4};
test_label[4702] = '{32'h42bb37aa};
test_output[4702] = '{32'h3f90f57e};
/*############ DEBUG ############
test_input[37616:37623] = '{-70.6598883096, 94.3522663162, -58.0221320827, 93.6087206782, -70.7925708323, -87.6742681029, -3.25544833346, 16.6030036416};
test_label[4702] = '{93.6087206782};
test_output[4702] = '{1.13249188308};
############ END DEBUG ############*/
test_input[37624:37631] = '{32'h4213cba1, 32'hc1d5a881, 32'hc22e2439, 32'hc1cf3220, 32'h428a94d8, 32'h422cc472, 32'hc1cf1d63, 32'hc26608e8};
test_label[4703] = '{32'hc22e2439};
test_output[4703] = '{32'h42e1a6f4};
/*############ DEBUG ############
test_input[37624:37631] = '{36.948855792, -26.7072772367, -43.5353750424, -25.8994753604, 69.2907086779, 43.19184209, -25.8893499348, -57.5086970151};
test_label[4703] = '{-43.5353750424};
test_output[4703] = '{112.82608372};
############ END DEBUG ############*/
test_input[37632:37639] = '{32'h40f25c27, 32'h42b62a63, 32'h429221f5, 32'hc295c9ac, 32'h4270bffc, 32'h41940beb, 32'h4250de9c, 32'h424ebe96};
test_label[4704] = '{32'h40f25c27};
test_output[4704] = '{32'h42a704a1};
/*############ DEBUG ############
test_input[37632:37639] = '{7.57374914624, 91.0827881373, 73.0663247586, -74.8938912117, 60.1874863542, 18.5058202179, 52.2173913097, 51.6861171893};
test_label[4704] = '{7.57374914624};
test_output[4704] = '{83.509039006};
############ END DEBUG ############*/
test_input[37640:37647] = '{32'hc1447a63, 32'hc2140415, 32'h42b0f342, 32'hc2844830, 32'h40d4abd6, 32'hc29f1c90, 32'hc2bbaae0, 32'hc284c70d};
test_label[4705] = '{32'hc2bbaae0};
test_output[4705] = '{32'h43364f11};
/*############ DEBUG ############
test_input[37640:37647] = '{-12.2798791853, -37.0039863202, 88.4751109875, -66.1409897972, 6.64597587146, -79.5557881819, -93.8337364331, -66.3887740394};
test_label[4705] = '{-93.8337364331};
test_output[4705] = '{182.308847421};
############ END DEBUG ############*/
test_input[37648:37655] = '{32'hc28509d0, 32'hc17a669d, 32'h4290ccf6, 32'hc26288ea, 32'h41a369ef, 32'h426d135b, 32'h42b91836, 32'h41bdad48};
test_label[4706] = '{32'h41a369ef};
test_output[4706] = '{32'h42903dba};
/*############ DEBUG ############
test_input[37648:37655] = '{-66.5191677254, -15.6500522833, 72.4003172592, -56.6337041246, 20.4267260809, 59.2689032174, 92.5472857467, 23.7096106469};
test_label[4706] = '{20.4267260809};
test_output[4706] = '{72.1205596676};
############ END DEBUG ############*/
test_input[37656:37663] = '{32'hc2c1779d, 32'hc1995d29, 32'h424cfd61, 32'hc284ee97, 32'hc2822ecf, 32'h41efa425, 32'h42b4e66e, 32'hc0b752a5};
test_label[4707] = '{32'h42b4e66e};
test_output[4707] = '{32'h80000000};
/*############ DEBUG ############
test_input[37656:37663] = '{-96.7336209099, -19.1704880023, 51.2474396636, -66.465995974, -65.0914241727, 29.9551485497, 90.4500609076, -5.72883845207};
test_label[4707] = '{90.4500609076};
test_output[4707] = '{-0.0};
############ END DEBUG ############*/
test_input[37664:37671] = '{32'h42be931f, 32'hc2c58ddc, 32'h418bf8a4, 32'hc2350474, 32'hc14b85ef, 32'h40cc9c48, 32'h42c023bc, 32'h4291f3fa};
test_label[4708] = '{32'hc2350474};
test_output[4708] = '{32'h430db362};
/*############ DEBUG ############
test_input[37664:37671] = '{95.2873477638, -98.7770722751, 17.4964063652, -45.2543492485, -12.7201985481, 6.39407709627, 96.0697948167, 72.9765200532};
test_label[4708] = '{-45.2543492485};
test_output[4708] = '{141.700719619};
############ END DEBUG ############*/
test_input[37672:37679] = '{32'h422d25a0, 32'hc268b0a1, 32'h427ae49d, 32'h41a2b166, 32'hc2529fba, 32'hc1aa9743, 32'hc0d52727, 32'hc1f23e5f};
test_label[4709] = '{32'hc2529fba};
test_output[4709] = '{32'h42e6c22b};
/*############ DEBUG ############
test_input[37672:37679] = '{43.2867418794, -58.1724874024, 62.7232541583, 20.3366194946, -52.6559815444, -21.3238577867, -6.66102942505, -30.2804542562};
test_label[4709] = '{-52.6559815444};
test_output[4709] = '{115.379235706};
############ END DEBUG ############*/
test_input[37680:37687] = '{32'hc1bfcd5e, 32'h425719a0, 32'hc29eaa2d, 32'hc22890b0, 32'hc29f6dc9, 32'h418c5e03, 32'h416c3903, 32'h418ed612};
test_label[4710] = '{32'hc1bfcd5e};
test_output[4710] = '{32'h429b8027};
/*############ DEBUG ############
test_input[37680:37687] = '{-23.9752770226, 53.7750225437, -79.3323708944, -42.1412963408, -79.7144217668, 17.5459050165, 14.7639184244, 17.8545259431};
test_label[4710] = '{-23.9752770226};
test_output[4710] = '{77.7502995663};
############ END DEBUG ############*/
test_input[37688:37695] = '{32'hc06609b4, 32'hc2a05767, 32'hc26fb1c2, 32'hc2007be3, 32'h4239ad13, 32'h42a70d6b, 32'hc1ed4d0a, 32'hc2a357a3};
test_label[4711] = '{32'h4239ad13};
test_output[4711] = '{32'h42146dc3};
/*############ DEBUG ############
test_input[37688:37695] = '{-3.59434221014, -80.1707056321, -59.9235922572, -32.1209842207, 46.4190196715, 83.5262071611, -29.6626175295, -81.6711677371};
test_label[4711] = '{46.4190196715};
test_output[4711] = '{37.1071874895};
############ END DEBUG ############*/
test_input[37696:37703] = '{32'h42a88368, 32'h42b1a773, 32'hc2bed317, 32'hc253b5b0, 32'hc249dafd, 32'hc1e4a993, 32'hc2b6fbd6, 32'hc22bce01};
test_label[4712] = '{32'hc2b6fbd6};
test_output[4712] = '{32'h43345448};
/*############ DEBUG ############
test_input[37696:37703] = '{84.2566501346, 88.827052023, -95.4122813856, -52.9274301949, -50.4638549321, -28.582799552, -91.4918694159, -42.9511742966};
test_label[4712] = '{-91.4918694159};
test_output[4712] = '{180.329222003};
############ END DEBUG ############*/
test_input[37704:37711] = '{32'h41a3ed3b, 32'hc2a9942e, 32'hc1e202ff, 32'h41ca9ef9, 32'h4294f99d, 32'hc21d9920, 32'hc2492fb4, 32'h42bea2f8};
test_label[4713] = '{32'hc2a9942e};
test_output[4713] = '{32'h43341b93};
/*############ DEBUG ############
test_input[37704:37711] = '{20.4908346549, -84.7894163705, -28.2514624592, 25.3276227063, 74.4875287641, -39.3995378616, -50.2965843968, 95.3183008268};
test_label[4713] = '{-84.7894163705};
test_output[4713] = '{180.107717198};
############ END DEBUG ############*/
test_input[37712:37719] = '{32'h42b0e7c6, 32'hc1ef9aa9, 32'h41e55e32, 32'hc0e47653, 32'hc293b508, 32'hc2673c4d, 32'h41139356, 32'h42b80c4d};
test_label[4714] = '{32'h42b80c4d};
test_output[4714] = '{32'h3ce329f1};
/*############ DEBUG ############
test_input[37712:37719] = '{88.4526827166, -29.9505177716, 28.6709936767, -7.13944403687, -73.8535788053, -57.8088871519, 9.2234703009, 92.0240275236};
test_label[4714] = '{92.0240275236};
test_output[4714] = '{0.0277299609695};
############ END DEBUG ############*/
test_input[37720:37727] = '{32'hc2a41a50, 32'hc293496a, 32'hc2b90216, 32'hc2655894, 32'hc2b68b49, 32'hc010aebb, 32'h4204023c, 32'h429f00d0};
test_label[4715] = '{32'hc2655894};
test_output[4715] = '{32'h4308d68d};
/*############ DEBUG ############
test_input[37720:37727] = '{-82.0513933871, -73.6433902852, -92.5040726994, -57.3365028227, -91.2720443431, -2.26066475247, 33.0021818422, 79.5015832121};
test_label[4715] = '{-57.3365028227};
test_output[4715] = '{136.838086035};
############ END DEBUG ############*/
test_input[37728:37735] = '{32'h42561ba9, 32'hc2363b05, 32'h42566d4d, 32'h40499be4, 32'h41ec2dee, 32'h41a9e218, 32'hc175ffc0, 32'hc20cd4a7};
test_label[4716] = '{32'hc20cd4a7};
test_output[4716] = '{32'h42b2efdd};
/*############ DEBUG ############
test_input[37728:37735] = '{53.5270130131, -45.5576360723, 53.6067387369, 3.15013981684, 29.5224272711, 21.2353975555, -15.3749389269, -35.2076683994};
test_label[4716] = '{-35.2076683994};
test_output[4716] = '{89.4684857686};
############ END DEBUG ############*/
test_input[37736:37743] = '{32'h42357682, 32'h41d5eff8, 32'hc1bd946a, 32'h42c58a7f, 32'h426df1a1, 32'hc2b4df73, 32'h429819da, 32'hc214fddc};
test_label[4717] = '{32'h426df1a1};
test_output[4717] = '{32'h421d235d};
/*############ DEBUG ############
test_input[37736:37743] = '{45.3657312453, 26.7421728788, -23.6974677132, 98.7705009978, 59.485964823, -90.4364218327, 76.0504905586, -37.2479111391};
test_label[4717] = '{59.485964823};
test_output[4717] = '{39.284536175};
############ END DEBUG ############*/
test_input[37744:37751] = '{32'hc26745e1, 32'h3f84d75b, 32'hc18b8bf2, 32'hc2b95667, 32'hc2a43a51, 32'hc2b7714c, 32'hc1e36121, 32'h42b4945e};
test_label[4718] = '{32'hc2b7714c};
test_output[4718] = '{32'h433602d5};
/*############ DEBUG ############
test_input[37744:37751] = '{-57.818239518, 1.03782213976, -17.4433321363, -92.6687522456, -82.1138984374, -91.721280595, -28.4224267293, 90.2897767231};
test_label[4718] = '{-91.721280595};
test_output[4718] = '{182.011057318};
############ END DEBUG ############*/
test_input[37752:37759] = '{32'hc2443120, 32'h42ad31d1, 32'hc1edb418, 32'hc24184ee, 32'hc1bdc937, 32'hc204a024, 32'hc196ac17, 32'h42a663c4};
test_label[4719] = '{32'hc204a024};
test_output[4719] = '{32'h42ef92a7};
/*############ DEBUG ############
test_input[37752:37759] = '{-49.0479751675, 86.597294739, -29.7129355852, -48.3798141127, -23.723250082, -33.1563880954, -18.8340276887, 83.1948522369};
test_label[4719] = '{-33.1563880954};
test_output[4719] = '{119.786432516};
############ END DEBUG ############*/
test_input[37760:37767] = '{32'hc1d5501d, 32'h4120d788, 32'hc0cf840f, 32'hc13c8d98, 32'h4215cc3d, 32'hc260ee99, 32'hc1ca2809, 32'h428b6a7b};
test_label[4720] = '{32'h4215cc3d};
test_output[4720] = '{32'h420108ba};
/*############ DEBUG ############
test_input[37760:37767] = '{-26.6641170281, 10.0526198086, -6.48487042096, -11.7845686949, 37.4494507495, -56.2330045854, -25.2695479749, 69.7079733833};
test_label[4720] = '{37.4494507495};
test_output[4720] = '{32.2585226338};
############ END DEBUG ############*/
test_input[37768:37775] = '{32'h42631f1c, 32'hc2c4645b, 32'hc207483d, 32'h41db873b, 32'h4180a3da, 32'hc1968548, 32'h422c181b, 32'hc2c41837};
test_label[4721] = '{32'h4180a3da};
test_output[4721] = '{32'h4222cd2f};
/*############ DEBUG ############
test_input[37768:37775] = '{56.7803816733, -98.1960040732, -33.8205448423, 27.4410309214, 16.0800064604, -18.8150780748, 43.0235393556, -98.0472909055};
test_label[4721] = '{16.0800064604};
test_output[4721] = '{40.7003762733};
############ END DEBUG ############*/
test_input[37776:37783] = '{32'h41b32a1a, 32'hc2482bff, 32'h42ba6776, 32'h4293af0b, 32'h42c34380, 32'h424605f2, 32'hc14d98f4, 32'hc24a70ba};
test_label[4722] = '{32'hc2482bff};
test_output[4722] = '{32'h4313afc8};
/*############ DEBUG ############
test_input[37776:37783] = '{22.3955574328, -50.0429653793, 93.2020693141, 73.8418808062, 97.6318387798, 49.5058063254, -12.8498425313, -50.6100840335};
test_label[4722] = '{-50.0429653793};
test_output[4722] = '{147.686650945};
############ END DEBUG ############*/
test_input[37784:37791] = '{32'hc19e6439, 32'hc260d6e2, 32'hc13c9878, 32'h42c2c4b2, 32'h42b51462, 32'h423404e2, 32'hc2395477, 32'hc1ea3d51};
test_label[4723] = '{32'hc2395477};
test_output[4723] = '{32'h430fb7bd};
/*############ DEBUG ############
test_input[37784:37791] = '{-19.7989377906, -56.2098447505, -11.7872240177, 97.3841714919, 90.5398127627, 45.0047675673, -46.3324858485, -29.2799387378};
test_label[4723] = '{-46.3324858485};
test_output[4723] = '{143.717722222};
############ END DEBUG ############*/
test_input[37792:37799] = '{32'hc1941fd4, 32'hc27ef629, 32'h4137b6f7, 32'h41c22f93, 32'h4126c346, 32'h42568e78, 32'hc2502526, 32'h42ad6483};
test_label[4724] = '{32'h42568e78};
test_output[4724] = '{32'h42043a8f};
/*############ DEBUG ############
test_input[37792:37799] = '{-18.5155417498, -63.7403923376, 11.4821690719, 24.2732290433, 10.4226738209, 53.6391279261, -52.0362783023, 86.6963149871};
test_label[4724] = '{53.6391279261};
test_output[4724] = '{33.057187061};
############ END DEBUG ############*/
test_input[37800:37807] = '{32'h42a546e0, 32'h427c9cfd, 32'hc2566386, 32'h42896763, 32'hc20b68b5, 32'h41c539ab, 32'hc2ace8c1, 32'hc24715f6};
test_label[4725] = '{32'h41c539ab};
test_output[4725] = '{32'h4267f0eb};
/*############ DEBUG ############
test_input[37800:37807] = '{82.6384279801, 63.1533097292, -53.5971918552, 68.7019273364, -34.852252138, 24.6531590549, -86.4545941372, -49.7714469795};
test_label[4725] = '{24.6531590549};
test_output[4725] = '{57.9852698147};
############ END DEBUG ############*/
test_input[37808:37815] = '{32'hc2c041da, 32'h4252faee, 32'h42a21c4c, 32'h4229e5a4, 32'hc28be43f, 32'hc0f94919, 32'h41d02850, 32'h40385793};
test_label[4726] = '{32'h40385793};
test_output[4726] = '{32'h429c598f};
/*############ DEBUG ############
test_input[37808:37815] = '{-96.1286134676, 52.7450468642, 81.0552671686, 42.4742589681, -69.9457912074, -7.79017318964, 26.0196839234, 2.88034506601};
test_label[4726] = '{2.88034506601};
test_output[4726] = '{78.1749221026};
############ END DEBUG ############*/
test_input[37816:37823] = '{32'hc1c42cb2, 32'h4286cb8d, 32'hc1d2a61d, 32'h42b180e4, 32'hc250f769, 32'h4294d51d, 32'hc293052c, 32'hc1253108};
test_label[4727] = '{32'h4294d51d};
test_output[4727] = '{32'h41655e38};
/*############ DEBUG ############
test_input[37816:37823] = '{-24.52182354, 67.3975579286, -26.3311101357, 88.751736297, -52.2416097391, 74.4162338261, -73.5101042706, -10.3244707305};
test_label[4727] = '{74.4162338261};
test_output[4727] = '{14.3355030659};
############ END DEBUG ############*/
test_input[37824:37831] = '{32'hc19ba9ce, 32'hc26895e1, 32'h42332e49, 32'hc23e28e7, 32'h4224dd52, 32'h42ac5246, 32'h4253de05, 32'h4272ba38};
test_label[4728] = '{32'h42332e49};
test_output[4728] = '{32'h42257644};
/*############ DEBUG ############
test_input[37824:37831] = '{-19.4579133558, -58.1463654482, 44.7951988121, -47.5399430467, 41.2161331869, 86.1606933262, 52.9668170778, 60.6818544655};
test_label[4728] = '{44.7951988121};
test_output[4728] = '{41.3654945141};
############ END DEBUG ############*/
test_input[37832:37839] = '{32'h429c6489, 32'hc26dfd75, 32'hc298423e, 32'h42228fbe, 32'h4126b9e7, 32'hc23b9975, 32'h41c5287d, 32'h420ebb44};
test_label[4729] = '{32'h429c6489};
test_output[4729] = '{32'h80000000};
/*############ DEBUG ############
test_input[37832:37839] = '{78.1963564749, -59.4975154423, -76.1293761083, 40.6403726107, 10.4203860501, -46.8998585541, 24.6447692738, 35.6828750504};
test_label[4729] = '{78.1963564749};
test_output[4729] = '{-0.0};
############ END DEBUG ############*/
test_input[37840:37847] = '{32'hc18b62b4, 32'hc280d3fc, 32'hc2307276, 32'hc28dfcc9, 32'h42a79c34, 32'hc20562bb, 32'h41897180, 32'h42b26f69};
test_label[4730] = '{32'h41897180};
test_output[4730] = '{32'h42901550};
/*############ DEBUG ############
test_input[37840:37847] = '{-17.4231954383, -64.4140346405, -44.1117770751, -70.9937185834, 83.8050810143, -33.3464173629, 17.1804207944, 89.217598615};
test_label[4730] = '{17.1804207944};
test_output[4730] = '{72.041628299};
############ END DEBUG ############*/
test_input[37848:37855] = '{32'hc2167496, 32'h42bd4605, 32'h42b7fe05, 32'hbed6544e, 32'h42951d57, 32'h4174aa16, 32'h41ec34d0, 32'h42976575};
test_label[4731] = '{32'hbed6544e};
test_output[4731] = '{32'h42be3f9f};
/*############ DEBUG ############
test_input[37848:37855] = '{-37.6138534949, 94.636758089, 91.9961340167, -0.418611945538, 74.5573074576, 15.2915246546, 29.525786899, 75.6981593645};
test_label[4731] = '{-0.418611945538};
test_output[4731] = '{95.1242585401};
############ END DEBUG ############*/
test_input[37856:37863] = '{32'h42a09288, 32'h42a4d2e3, 32'h41c5d2e4, 32'hc120c9ca, 32'hc1872424, 32'hc2030965, 32'h42b53a7c, 32'h429d96c5};
test_label[4732] = '{32'h41c5d2e4};
test_output[4732] = '{32'h4283c5ed};
/*############ DEBUG ############
test_input[37856:37863] = '{80.2861911836, 82.4118866975, 24.7279730192, -10.0492652307, -16.8926460959, -32.7591736387, 90.6142302719, 78.7944727565};
test_label[4732] = '{24.7279730192};
test_output[4732] = '{65.886571275};
############ END DEBUG ############*/
test_input[37864:37871] = '{32'hc2b54b58, 32'h41ee88e6, 32'h41a2438e, 32'hc274587c, 32'h41503f4c, 32'hc258b8ff, 32'hc254d762, 32'h3fbb7563};
test_label[4733] = '{32'h41ee88e6};
test_output[4733] = '{32'h3897d992};
/*############ DEBUG ############
test_input[37864:37871] = '{-90.6471569893, 29.81684549, 20.2829857603, -61.0864106982, 13.0154533722, -54.1806598168, -53.2103339297, 1.46451988484};
test_label[4733] = '{29.81684549};
test_output[4733] = '{7.24076690125e-05};
############ END DEBUG ############*/
test_input[37872:37879] = '{32'h411db319, 32'hc26ecc4a, 32'h4292c8bd, 32'h4109d996, 32'hc28a7d5c, 32'h42baa47d, 32'h42aeeb0f, 32'h41ecaaa1};
test_label[4734] = '{32'h41ecaaa1};
test_output[4734] = '{32'h427ef693};
/*############ DEBUG ############
test_input[37872:37879] = '{9.85622457323, -59.6994993935, 73.392065201, 8.61562113499, -69.244839102, 93.3212677978, 87.4590955927, 29.58331411};
test_label[4734] = '{29.58331411};
test_output[4734] = '{63.7407947074};
############ END DEBUG ############*/
test_input[37880:37887] = '{32'hc1f7f758, 32'hc2a60a0e, 32'h41b3ae7f, 32'h42700240, 32'hc2818c10, 32'h42ae7e97, 32'hc2b631a7, 32'hc0f46ef5};
test_label[4735] = '{32'hc2a60a0e};
test_output[4735] = '{32'h432a4452};
/*############ DEBUG ############
test_input[37880:37887] = '{-30.9957735731, -83.0196380527, 22.4602022577, 60.0021981898, -64.7735597776, 87.2472432189, -91.0969740144, -7.63854462244};
test_label[4735] = '{-83.0196380527};
test_output[4735] = '{170.266881272};
############ END DEBUG ############*/
test_input[37888:37895] = '{32'h4283099e, 32'h427a4f16, 32'h421cf8ad, 32'h42c59553, 32'h4166ee6e, 32'hc217c7d0, 32'hc17ce662, 32'h42266ce4};
test_label[4736] = '{32'h4283099e};
test_output[4736] = '{32'h4205176a};
/*############ DEBUG ############
test_input[37888:37895] = '{65.5187816824, 62.5772324872, 39.2428488463, 98.7916463117, 14.433210319, -37.9451301835, -15.8062457994, 41.60633681};
test_label[4736] = '{65.5187816824};
test_output[4736] = '{33.2728646293};
############ END DEBUG ############*/
test_input[37896:37903] = '{32'h42867a1a, 32'hc2b5157f, 32'h429ce6ae, 32'hc290dfed, 32'h42b964aa, 32'hc2b09446, 32'hc2b2fe50, 32'hc28e630e};
test_label[4737] = '{32'h42867a1a};
test_output[4737] = '{32'h41cbaa43};
/*############ DEBUG ############
test_input[37896:37903] = '{67.2384760032, -90.5419839387, 78.4505460682, -72.4373521457, 92.6966113198, -88.2895945053, -89.4967055112, -71.1934672911};
test_label[4737] = '{67.2384760032};
test_output[4737] = '{25.4581359668};
############ END DEBUG ############*/
test_input[37904:37911] = '{32'hc12bfda9, 32'hc2075647, 32'h422b9168, 32'hc2a0c840, 32'h42c56994, 32'h401d7dbd, 32'h3d2f472c, 32'h42bb9fd6};
test_label[4738] = '{32'h42bb9fd6};
test_output[4738] = '{32'h409cd906};
/*############ DEBUG ############
test_input[37904:37911] = '{-10.7494288279, -33.8342562825, 42.8919984911, -80.3911168179, 98.706208228, 2.46079936962, 0.0427924842147, 93.8121791823};
test_label[4738] = '{93.8121791823};
test_output[4738] = '{4.90149230549};
############ END DEBUG ############*/
test_input[37912:37919] = '{32'hc0877d69, 32'hc105925b, 32'h42b5563f, 32'hc2c2a695, 32'hc25cc964, 32'h409cad53, 32'h427178a2, 32'hc198d13e};
test_label[4739] = '{32'hc105925b};
test_output[4739] = '{32'h42c6088a};
/*############ DEBUG ############
test_input[37912:37919] = '{-4.23405890062, -8.34823145592, 90.6684464283, -97.3253520191, -55.1966712598, 4.89615759251, 60.3678049132, -19.1021699723};
test_label[4739] = '{-8.34823145592};
test_output[4739] = '{99.0166778843};
############ END DEBUG ############*/
test_input[37920:37927] = '{32'hc26c3564, 32'hc1ebbc31, 32'h41864e4d, 32'h41fa064a, 32'hc2b01b5b, 32'hc11523e8, 32'h4262c8eb, 32'h42c7c24e};
test_label[4740] = '{32'h42c7c24e};
test_output[4740] = '{32'h80000000};
/*############ DEBUG ############
test_input[37920:37927] = '{-59.0521385773, -29.4668894409, 16.7882332441, 31.2530709707, -88.0534253714, -9.32126571664, 56.6962084387, 99.8794976439};
test_label[4740] = '{99.8794976439};
test_output[4740] = '{-0.0};
############ END DEBUG ############*/
test_input[37928:37935] = '{32'h423ae19b, 32'hc298f579, 32'hc2af71b0, 32'hc23c5084, 32'hc130322e, 32'hc18e9535, 32'hc1ae931e, 32'h42677106};
test_label[4741] = '{32'h423ae19b};
test_output[4741] = '{32'h41323dbe};
/*############ DEBUG ############
test_input[37928:37935] = '{46.7203168922, -76.479441871, -87.7220451448, -47.0786285492, -11.0122510959, -17.822854525, -21.8218352824, 57.8603759196};
test_label[4741] = '{46.7203168922};
test_output[4741] = '{11.1400735463};
############ END DEBUG ############*/
test_input[37936:37943] = '{32'hc268ecbf, 32'hc0843d18, 32'hc28c774d, 32'h4248cd9d, 32'h410f9f70, 32'hc28cfd86, 32'h428cc5cf, 32'hbf905eb2};
test_label[4742] = '{32'hc28c774d};
test_output[4742] = '{32'h430c9e8e};
/*############ DEBUG ############
test_input[37936:37943] = '{-58.2311991912, -4.13245773813, -70.2330094507, 50.2007948629, 8.97642507667, -70.495166685, 70.386343057, -1.12788990009};
test_label[4742] = '{-70.2330094507};
test_output[4742] = '{140.619352509};
############ END DEBUG ############*/
test_input[37944:37951] = '{32'hc2a4419f, 32'hc063481c, 32'h4243d90d, 32'hc260c85f, 32'hc22ca1bf, 32'h424fd30c, 32'h429b9ec8, 32'hc2b299d3};
test_label[4743] = '{32'h4243d90d};
test_output[4743] = '{32'h41e6c908};
/*############ DEBUG ############
test_input[37944:37951] = '{-82.1281669664, -3.55127622405, 48.9619634275, -56.1956761597, -43.157955277, 51.9561004251, 77.8101231929, -89.3004372943};
test_label[4743] = '{48.9619634275};
test_output[4743] = '{28.8481597654};
############ END DEBUG ############*/
test_input[37952:37959] = '{32'hc210ed89, 32'hc1fbf7f4, 32'hc297481c, 32'hc1c7092a, 32'hc2a2c810, 32'h421fb2e6, 32'h41eda35d, 32'hc2b07cc9};
test_label[4744] = '{32'hc297481c};
test_output[4744] = '{32'h42e72194};
/*############ DEBUG ############
test_input[37952:37959] = '{-36.2319673835, -31.4960705353, -75.6408357236, -24.879475026, -81.3907469853, 39.9247068093, 29.7047673392, -88.2437175568};
test_label[4744] = '{-75.6408357236};
test_output[4744] = '{115.565578969};
############ END DEBUG ############*/
test_input[37960:37967] = '{32'h42a633d5, 32'hc0baf590, 32'h4211a3e8, 32'hc2048af1, 32'hc2accff9, 32'hc28d342f, 32'hc231b36f, 32'h42c63594};
test_label[4745] = '{32'hc0baf590};
test_output[4745] = '{32'h42d1e4ed};
/*############ DEBUG ############
test_input[37960:37967] = '{83.101234337, -5.84247584784, 36.4100664931, -33.1356857795, -86.4061962332, -70.601918702, -44.4252297783, 99.1046415473};
test_label[4745] = '{-5.84247584784};
test_output[4745] = '{104.947117507};
############ END DEBUG ############*/
test_input[37968:37975] = '{32'h415203f0, 32'hc257c767, 32'hc2554c34, 32'h425539b7, 32'h41a341eb, 32'h408e844c, 32'hc1af708c, 32'hc24eab4b};
test_label[4746] = '{32'h425539b7};
test_output[4746] = '{32'h27b80000};
/*############ DEBUG ############
test_input[37968:37975] = '{13.125961191, -53.9447269473, -53.3244170173, 53.3063608439, 20.4071858981, 4.45364960907, -21.9299540323, -51.6672796888};
test_label[4746] = '{53.3063608439};
test_output[4746] = '{5.10702591328e-15};
############ END DEBUG ############*/
test_input[37976:37983] = '{32'h42b6cf17, 32'h42bade8c, 32'h42b72fc2, 32'hc2484e10, 32'h42094891, 32'h425e23f1, 32'h42ae05c9, 32'hc20cbc47};
test_label[4747] = '{32'h42ae05c9};
test_output[4747] = '{32'h40d5bbe3};
/*############ DEBUG ############
test_input[37976:37983] = '{91.4044714036, 93.434658406, 91.5932786484, -50.0762329883, 34.3208648583, 55.535098663, 87.0113024056, -35.1838650815};
test_label[4747] = '{87.0113024056};
test_output[4747] = '{6.67918558384};
############ END DEBUG ############*/
test_input[37984:37991] = '{32'h416b8a1f, 32'h427eba58, 32'h41ca4d92, 32'hc2bc5140, 32'hc1900fb7, 32'h426487c1, 32'hc23745f8, 32'h4222cac7};
test_label[4748] = '{32'hc2bc5140};
test_output[4748] = '{32'h431dd794};
/*############ DEBUG ############
test_input[37984:37991] = '{14.7212213446, 63.6819750192, 25.287875892, -94.158692608, -18.0076733583, 57.1325705809, -45.8183278947, 40.6980239041};
test_label[4748] = '{-94.158692608};
test_output[4748] = '{157.842097572};
############ END DEBUG ############*/
test_input[37992:37999] = '{32'h42360066, 32'h42b9633f, 32'hc2a01e19, 32'hc253a696, 32'hc196861c, 32'h428723f9, 32'h41aab812, 32'hc22446cd};
test_label[4749] = '{32'h428723f9};
test_output[4749] = '{32'h41c8fd19};
/*############ DEBUG ############
test_input[37992:37999] = '{45.500390617, 92.6938414145, -80.0587841741, -52.9126830334, -18.8154833166, 67.5702594369, 21.3398778815, -41.0691420135};
test_label[4749] = '{67.5702594369};
test_output[4749] = '{25.1235819775};
############ END DEBUG ############*/
test_input[38000:38007] = '{32'hc26d1c4b, 32'hc16da912, 32'hc2832841, 32'h4108d49c, 32'hc2922300, 32'hc2bf0ddd, 32'h4285699b, 32'hc2a56977};
test_label[4750] = '{32'hc2832841};
test_output[4750] = '{32'h430448ee};
/*############ DEBUG ############
test_input[38000:38007] = '{-59.2776286225, -14.853776679, -65.5786238452, 8.55190641696, -73.0683599305, -95.5270803441, 66.7062638046, -82.705982956};
test_label[4750] = '{-65.5786238452};
test_output[4750] = '{132.28488765};
############ END DEBUG ############*/
test_input[38008:38015] = '{32'hc2505d49, 32'hc23d7424, 32'hc28dd006, 32'h4232ed28, 32'h4299d961, 32'h4162cceb, 32'hc2255025, 32'hc2a73fa4};
test_label[4751] = '{32'hc28dd006};
test_output[4751] = '{32'h4313d4b3};
/*############ DEBUG ############
test_input[38008:38015] = '{-52.0910995085, -47.3634180384, -70.906292807, 44.7315963275, 76.9245710159, 14.1750291993, -41.3282665861, -83.6242980254};
test_label[4751] = '{-70.906292807};
test_output[4751] = '{147.830863823};
############ END DEBUG ############*/
test_input[38016:38023] = '{32'h424b9e21, 32'hc21e9a17, 32'hc21534f4, 32'h42b95270, 32'hc21c6167, 32'h416cb78b, 32'h41934bbf, 32'h4184623a};
test_label[4752] = '{32'h41934bbf};
test_output[4752] = '{32'h42947f80};
/*############ DEBUG ############
test_input[38016:38023] = '{50.9044240718, -39.6504785515, -37.3017120086, 92.6610079379, -39.0951208971, 14.7948098279, 18.4119852911, 16.5479619845};
test_label[4752] = '{18.4119852911};
test_output[4752] = '{74.2490226469};
############ END DEBUG ############*/
test_input[38024:38031] = '{32'hc25e6a14, 32'h42784cd8, 32'hc22d69f6, 32'hc23beb6c, 32'h42a9caf7, 32'hc26ea796, 32'hc220cb4f, 32'h41c30c31};
test_label[4753] = '{32'h42a9caf7};
test_output[4753] = '{32'h2f06e5b0};
/*############ DEBUG ############
test_input[38024:38031] = '{-55.6035915887, 62.0750445331, -43.3534785963, -46.9799049562, 84.8964187666, -59.6636575661, -40.1985430037, 24.3809526543};
test_label[4753] = '{84.8964187666};
test_output[4753] = '{1.22688303968e-10};
############ END DEBUG ############*/
test_input[38032:38039] = '{32'hc29a2d9f, 32'hc2bbc2ac, 32'hc2881f89, 32'h428f29af, 32'hc2b48d05, 32'h420020f6, 32'hc2362ca5, 32'h42583a6e};
test_label[4754] = '{32'hc2b48d05};
test_output[4754] = '{32'h4321db5a};
/*############ DEBUG ############
test_input[38032:38039] = '{-77.0891042219, -93.8802150802, -68.0615935775, 71.5814153716, -90.2754251048, 32.0321866027, -45.5435983389, 54.057060641};
test_label[4754] = '{-90.2754251048};
test_output[4754] = '{161.856840501};
############ END DEBUG ############*/
test_input[38040:38047] = '{32'h42643c7c, 32'h42ac8b38, 32'hc2aef283, 32'hc251b68e, 32'h426a6428, 32'hc12483cc, 32'hc2c4697e, 32'hbfc9f715};
test_label[4755] = '{32'h426a6428};
test_output[4755] = '{32'h41dd648f};
/*############ DEBUG ############
test_input[38040:38047] = '{57.0590650777, 86.2719083095, -87.4736551553, -52.4282765982, 58.597807757, -10.282177416, -98.2060417144, -1.57785279878};
test_label[4755] = '{58.597807757};
test_output[4755] = '{27.6741005525};
############ END DEBUG ############*/
test_input[38048:38055] = '{32'hc237f68f, 32'hc299e8a8, 32'hc2951459, 32'h426c858e, 32'hc202083e, 32'hc24bea53, 32'h4159830b, 32'h4293d990};
test_label[4756] = '{32'hc299e8a8};
test_output[4756] = '{32'h4316e11c};
/*############ DEBUG ############
test_input[38048:38055] = '{-45.9907782145, -76.9544053798, -74.5397440314, 59.1304238529, -32.5080480791, -50.9788335928, 13.5944929424, 73.9249233839};
test_label[4756] = '{-76.9544053798};
test_output[4756] = '{150.879329139};
############ END DEBUG ############*/
test_input[38056:38063] = '{32'hc292f14f, 32'hc1df3d9e, 32'hc2a8b506, 32'h41aee157, 32'h4276ddfe, 32'h42086fc0, 32'h4246e8de, 32'h42bfc891};
test_label[4757] = '{32'h41aee157};
test_output[4757] = '{32'h4294103b};
/*############ DEBUG ############
test_input[38056:38063] = '{-73.4713059966, -27.9050873678, -84.3535608259, 21.86003003, 61.7167908658, 34.1091295942, 49.7274090059, 95.8917306207};
test_label[4757] = '{21.86003003};
test_output[4757] = '{74.0317005908};
############ END DEBUG ############*/
test_input[38064:38071] = '{32'h42c5b9f9, 32'h429f47e0, 32'h415f7d2a, 32'hc1f67b06, 32'hc277383a, 32'h422aa189, 32'h422b8e60, 32'h42468963};
test_label[4758] = '{32'h42468963};
test_output[4758] = '{32'h4244ea8f};
/*############ DEBUG ############
test_input[38064:38071] = '{98.8632293174, 79.6403813911, 13.9680572945, -30.8100699225, -61.8049072265, 42.6577503343, 42.8890397453, 49.6341674593};
test_label[4758] = '{49.6341674593};
test_output[4758] = '{49.2290618625};
############ END DEBUG ############*/
test_input[38072:38079] = '{32'h42b2e756, 32'hc26d3089, 32'hc1dd5b5f, 32'hc2abf20c, 32'hc2ae7668, 32'hc21f7e5b, 32'h41ea65fe, 32'hc2b566ee};
test_label[4759] = '{32'hc21f7e5b};
test_output[4759] = '{32'h43015342};
/*############ DEBUG ############
test_input[38072:38079] = '{89.4518296417, -59.2973963125, -27.669614262, -85.9727440026, -87.2312648463, -39.8733954454, 29.2998017129, -90.7010310038};
test_label[4759] = '{-39.8733954454};
test_output[4759] = '{129.325225087};
############ END DEBUG ############*/
test_input[38080:38087] = '{32'hc28c5dc3, 32'hc2381098, 32'h4208783a, 32'h421d3b6d, 32'hc1b2bece, 32'h4143a645, 32'hc172d73b, 32'h42441618};
test_label[4760] = '{32'hc28c5dc3};
test_output[4760] = '{32'h42ee68d7};
/*############ DEBUG ############
test_input[38080:38087] = '{-70.1831266584, -46.0162044226, 34.1174083486, 39.3080326198, -22.3431671751, 12.2280932723, -15.1775461695, 49.0215769199};
test_label[4760] = '{-70.1831266584};
test_output[4760] = '{119.204764372};
############ END DEBUG ############*/
test_input[38088:38095] = '{32'hc23f37c6, 32'hc29b346a, 32'h42c47835, 32'hc26c09b0, 32'h42bbd708, 32'h420662fd, 32'hc1f12331, 32'h42a55fa4};
test_label[4761] = '{32'h42c47835};
test_output[4761] = '{32'h3c599815};
/*############ DEBUG ############
test_input[38088:38095] = '{-47.8044665145, -77.6023709927, 98.2347769478, -59.009461671, 93.9199822753, 33.5966665726, -30.1421840587, 82.6867978486};
test_label[4761] = '{98.2347769478};
test_output[4761] = '{0.0132808884188};
############ END DEBUG ############*/
test_input[38096:38103] = '{32'hbe0b0b40, 32'hc28a840d, 32'h42af5d25, 32'h42b3d84e, 32'h428502fb, 32'hc20d8502, 32'h42575adb, 32'hc196e4e0};
test_label[4762] = '{32'hc196e4e0};
test_output[4762] = '{32'h42d9c54a};
/*############ DEBUG ############
test_input[38096:38103] = '{-0.135785109412, -69.2579089377, 87.6819240955, 89.9224663253, 66.5058190488, -35.3798917767, 53.8387264355, -18.8617552281};
test_label[4762] = '{-18.8617552281};
test_output[4762] = '{108.885333773};
############ END DEBUG ############*/
test_input[38104:38111] = '{32'h4144b27d, 32'hc19ae055, 32'h42a2a6e8, 32'h414aa954, 32'hc1183bbe, 32'h42b2d6ba, 32'hc2009f55, 32'hc21a15b0};
test_label[4763] = '{32'hc1183bbe};
test_output[4763] = '{32'h42c5de5a};
/*############ DEBUG ############
test_input[38104:38111] = '{12.2935767087, -19.3595377175, 81.3259893414, 12.6663400413, -9.51458550473, 89.4193914487, -32.1555989815, -38.521177552};
test_label[4763] = '{-9.51458550473};
test_output[4763] = '{98.9342824552};
############ END DEBUG ############*/
test_input[38112:38119] = '{32'hc266dfa2, 32'hc1173712, 32'hc1e17166, 32'hc21d0309, 32'hc27919f0, 32'h4208ef0c, 32'hc18cab09, 32'h42b02d7a};
test_label[4764] = '{32'hc27919f0};
test_output[4764] = '{32'h43165d39};
/*############ DEBUG ############
test_input[38112:38119] = '{-57.718393259, -9.45094467777, -28.1803708292, -39.2529627446, -62.2753286615, 34.2334439052, -17.5835125127, 88.0888188514};
test_label[4764] = '{-62.2753286615};
test_output[4764] = '{150.364147513};
############ END DEBUG ############*/
test_input[38120:38127] = '{32'h423927f1, 32'hc28ce6c7, 32'h429d2fe6, 32'h425ae499, 32'h41a1929a, 32'h42728bc6, 32'hc1320026, 32'h41cbe2d6};
test_label[4765] = '{32'hc1320026};
test_output[4765] = '{32'h42b36fea};
/*############ DEBUG ############
test_input[38120:38127] = '{46.2890067383, -70.4507352854, 78.5935481574, 54.7232381164, 20.1965833287, 60.6364977656, -11.1250364699, 25.4857596419};
test_label[4765] = '{-11.1250364699};
test_output[4765] = '{89.7185846432};
############ END DEBUG ############*/
test_input[38128:38135] = '{32'h42b05dfa, 32'h42694daf, 32'hc28b71db, 32'hc29f5a14, 32'h42a6b472, 32'hc1eacd87, 32'h42b3c2ca, 32'h422eaa93};
test_label[4766] = '{32'h42b3c2ca};
test_output[4766] = '{32'h3e2d91a6};
/*############ DEBUG ############
test_input[38128:38135] = '{88.183549582, 58.3258614812, -69.7223755394, -79.6759315548, 83.3524313025, -29.3503554727, 89.8804451772, 43.6665765061};
test_label[4766] = '{89.8804451772};
test_output[4766] = '{0.169500918632};
############ END DEBUG ############*/
test_input[38136:38143] = '{32'hc1dc9386, 32'h40870dad, 32'h42b3db3f, 32'hc2a59e53, 32'h41c5f833, 32'h4224d2c0, 32'hc2559848, 32'h417cbbdd};
test_label[4767] = '{32'hc1dc9386};
test_output[4767] = '{32'h42eb0021};
/*############ DEBUG ############
test_input[38136:38143] = '{-27.5720323765, 4.2204193645, 89.928218552, -82.8092299481, 24.7461918951, 41.2058099139, -53.3987133245, 15.7958653062};
test_label[4767] = '{-27.5720323765};
test_output[4767] = '{117.500250928};
############ END DEBUG ############*/
test_input[38144:38151] = '{32'h4258481e, 32'h428bdd7f, 32'hc1c7f198, 32'hc2bd6122, 32'hc2138456, 32'h41da182b, 32'hc23420fe, 32'hc29f63ec};
test_label[4768] = '{32'hc1c7f198};
test_output[4768] = '{32'h42bdd9e5};
/*############ DEBUG ############
test_input[38144:38151] = '{54.07042571, 69.9326071398, -24.9929659287, -94.6897140616, -36.8792332671, 27.2618000622, -45.0322177666, -79.695159791};
test_label[4768] = '{-24.9929659287};
test_output[4768] = '{94.9255731976};
############ END DEBUG ############*/
test_input[38152:38159] = '{32'hc2be401c, 32'h42b620ab, 32'h42343de7, 32'hc117c5fe, 32'h41494227, 32'h4200f7c8, 32'hbfbbd5f0, 32'h42ad67f8};
test_label[4769] = '{32'hbfbbd5f0};
test_output[4769] = '{32'h42b91682};
/*############ DEBUG ############
test_input[38152:38159] = '{-95.125212161, 91.0638048592, 45.0604516664, -9.48583819121, 12.5786505479, 32.2419745814, -1.46746637279, 86.7030658472};
test_label[4769] = '{-1.46746637279};
test_output[4769] = '{92.5439593441};
############ END DEBUG ############*/
test_input[38160:38167] = '{32'hc1e9d022, 32'h40d08f5c, 32'hc19622bd, 32'hc2c138b5, 32'h42617982, 32'h422a4792, 32'hc2a66236, 32'h42b9289a};
test_label[4770] = '{32'h42617982};
test_output[4770] = '{32'h4210d7b3};
/*############ DEBUG ############
test_input[38160:38167] = '{-29.2266268389, 6.51749998769, -18.766962914, -96.6107585744, 56.3686589474, 42.569893159, -83.1918153679, 92.5793030131};
test_label[4770] = '{56.3686589474};
test_output[4770] = '{36.2106440657};
############ END DEBUG ############*/
test_input[38168:38175] = '{32'hc281ae42, 32'hc20fbaaa, 32'hc1f30684, 32'h3e48f5a0, 32'hc29b7ae9, 32'hc2459652, 32'h427454a9, 32'h4296d697};
test_label[4771] = '{32'hc281ae42};
test_output[4771] = '{32'h430c426d};
/*############ DEBUG ############
test_input[38168:38175] = '{-64.8403497135, -35.9322892695, -30.3781808159, 0.196249481072, -77.7400575337, -49.396796913, 61.0826742108, 75.4191199425};
test_label[4771] = '{-64.8403497135};
test_output[4771] = '{140.25947025};
############ END DEBUG ############*/
test_input[38176:38183] = '{32'hc211cdd2, 32'h40331d21, 32'hc28de889, 32'hc285f1b5, 32'hc2229481, 32'h4259cee3, 32'hc23c787a, 32'hc2c3480a};
test_label[4772] = '{32'h40331d21};
test_output[4772] = '{32'h424e9d11};
/*############ DEBUG ############
test_input[38176:38183] = '{-36.4509958508, 2.79865300171, -70.954172845, -66.972082101, -40.6450227214, 54.4520390346, -47.1176523579, -97.6406999119};
test_label[4772] = '{2.79865300171};
test_output[4772] = '{51.6533860329};
############ END DEBUG ############*/
test_input[38184:38191] = '{32'hc1809a6e, 32'h429cef6e, 32'h42b325c7, 32'h41e7bbcc, 32'hc293203e, 32'h429b8b44, 32'h427d01a9, 32'hc274bcf3};
test_label[4773] = '{32'hc1809a6e};
test_output[4773] = '{32'h42d34c66};
/*############ DEBUG ############
test_input[38184:38191] = '{-16.0754044329, 78.4676352391, 89.5737858231, 28.9666976983, -73.5629696964, 77.7719999854, 63.2516230649, -61.1845220841};
test_label[4773] = '{-16.0754044329};
test_output[4773] = '{105.649212767};
############ END DEBUG ############*/
test_input[38192:38199] = '{32'hc1c25064, 32'h42abaf36, 32'hc2ac7ee3, 32'h4269d0fc, 32'h42283742, 32'h42998de9, 32'h42bd9cd9, 32'hc247e386};
test_label[4774] = '{32'h42283742};
test_output[4774] = '{32'h42530291};
/*############ DEBUG ############
test_input[38192:38199] = '{-24.2892531406, 85.8422053488, -86.2478234471, 58.4540846845, 42.0539630539, 76.7771697254, 94.8063418214, -49.9721903626};
test_label[4774] = '{42.0539630539};
test_output[4774] = '{52.7525066902};
############ END DEBUG ############*/
test_input[38200:38207] = '{32'h42abf1bf, 32'hbf7e4dda, 32'hc16372f2, 32'hc2c10fd1, 32'hc23bbb21, 32'h429fc17c, 32'hc2ae25df, 32'h4204f192};
test_label[4775] = '{32'hc16372f2};
test_output[4775] = '{32'h42c86144};
/*############ DEBUG ############
test_input[38200:38207] = '{85.9721592171, -0.993375404275, -14.2155624186, -96.5308915762, -46.9327439384, 79.8779006274, -87.0739665486, 33.2359085192};
test_label[4775] = '{-14.2155624186};
test_output[4775] = '{100.189974877};
############ END DEBUG ############*/
test_input[38208:38215] = '{32'hc2ae3f1f, 32'h42b07ef4, 32'h42bc22a1, 32'h4298b670, 32'hc15fbb37, 32'hc29dec18, 32'hc2a99479, 32'h42b631ed};
test_label[4776] = '{32'h42b631ed};
test_output[4776] = '{32'h40417860};
/*############ DEBUG ############
test_input[38208:38215] = '{-87.1232818249, 88.2479579585, 94.067637258, 76.356322178, -13.9832070711, -78.9611241066, -84.7899879014, 91.0975092459};
test_label[4776] = '{91.0975092459};
test_output[4776] = '{3.0229721579};
############ END DEBUG ############*/
test_input[38216:38223] = '{32'hc293b47a, 32'hbf329202, 32'h42b8a9a3, 32'h40c7e659, 32'hc29043a5, 32'h41ee44af, 32'hc1b30934, 32'h42738a25};
test_label[4777] = '{32'h42738a25};
test_output[4777] = '{32'h41fb9242};
/*############ DEBUG ############
test_input[38216:38223] = '{-73.8524958579, -0.697540396208, 92.3313195183, 6.24686883007, -72.1321176569, 29.7835365717, -22.3794937496, 60.8849050885};
test_label[4777] = '{60.8849050885};
test_output[4777] = '{31.4464144298};
############ END DEBUG ############*/
test_input[38224:38231] = '{32'hc2b93b4c, 32'hc2289a52, 32'h41f7d89a, 32'h42650b49, 32'hc2a89831, 32'h426fb31c, 32'h407cad05, 32'h42b2a6fe};
test_label[4778] = '{32'h41f7d89a};
test_output[4778] = '{32'h426961ae};
/*############ DEBUG ############
test_input[38224:38231] = '{-92.6158107846, -42.1507049517, 30.9807632904, 57.2610196277, -84.2972503914, 59.9249106555, 3.94806034439, 89.3261551924};
test_label[4778] = '{30.9807632904};
test_output[4778] = '{58.345391902};
############ END DEBUG ############*/
test_input[38232:38239] = '{32'h423fac62, 32'h41af9fe5, 32'hc2c15212, 32'h425d17cc, 32'hc2860385, 32'h415636f7, 32'hc2c087a7, 32'h42af0e54};
test_label[4779] = '{32'hc2c15212};
test_output[4779] = '{32'h43383033};
/*############ DEBUG ############
test_input[38232:38239] = '{47.9183408313, 21.9530736249, -96.6602953346, 55.2732405552, -67.0068706708, 13.3884187034, -96.2649464883, 87.5279811324};
test_label[4779] = '{-96.6602953346};
test_output[4779] = '{184.188276467};
############ END DEBUG ############*/
test_input[38240:38247] = '{32'hc2b9a0a8, 32'h426feb3b, 32'h4299f81d, 32'h42a7f0be, 32'hc1e950ff, 32'h4245dc02, 32'h4202823e, 32'h420cf917};
test_label[4780] = '{32'h426feb3b};
test_output[4780] = '{32'h41bfee67};
/*############ DEBUG ############
test_input[38240:38247] = '{-92.8137855509, 59.979716679, 76.9845953454, 83.970198864, -29.1645495492, 49.4648507917, 32.6271880175, 35.2432529182};
test_label[4780] = '{59.979716679};
test_output[4780] = '{23.9914068622};
############ END DEBUG ############*/
test_input[38248:38255] = '{32'h40f80d42, 32'hc2b6c3d8, 32'hc28786a2, 32'h42145e2d, 32'h404452e5, 32'hc2114548, 32'h4226b81f, 32'h40db2d3d};
test_label[4781] = '{32'h404452e5};
test_output[4781] = '{32'h421a7d4f};
/*############ DEBUG ############
test_input[38248:38255] = '{7.75161855721, -91.3825058729, -67.7629580334, 37.0919666585, 3.06755941911, -36.3176582198, 41.6798072011, 6.84927214084};
test_label[4781] = '{3.06755941911};
test_output[4781] = '{38.6223711738};
############ END DEBUG ############*/
test_input[38256:38263] = '{32'hc26a86b2, 32'h42a48acd, 32'h42a819e4, 32'hc299556b, 32'hc29a2efd, 32'h4253eab3, 32'hc20f304e, 32'hc196cc4b};
test_label[4782] = '{32'hc299556b};
test_output[4782] = '{32'h4320df92};
/*############ DEBUG ############
test_input[38256:38263] = '{-58.6315381834, 82.2710976998, 84.0505674159, -76.6668341236, -77.0917707857, 52.9791984789, -35.7971710083, -18.849751702};
test_label[4782] = '{-76.6668341236};
test_output[4782] = '{160.873317173};
############ END DEBUG ############*/
test_input[38264:38271] = '{32'hc23d8abc, 32'h422cfa0b, 32'hc291f4a9, 32'hc2bec6cb, 32'h4283b51d, 32'hc2249f4b, 32'h42862b22, 32'h4283ef09};
test_label[4783] = '{32'h42862b22};
test_output[4783] = '{32'h3ef6c670};
/*############ DEBUG ############
test_input[38264:38271] = '{-47.385482953, 43.244181364, -72.9778536026, -95.388264042, 65.8537359932, -41.155557912, 67.0842423348, 65.9668665507};
test_label[4783] = '{67.0842423348};
test_output[4783] = '{0.481982694766};
############ END DEBUG ############*/
test_input[38272:38279] = '{32'h41b2f41b, 32'hc2956db9, 32'h428a2e99, 32'hc22b63b4, 32'hc13881ce, 32'hc286e88f, 32'h42bf23ab, 32'hc1ef98de};
test_label[4784] = '{32'hc286e88f};
test_output[4784] = '{32'h4323061d};
/*############ DEBUG ############
test_input[38272:38279] = '{22.3691925666, -74.7143042406, 69.0910109811, -42.8473677636, -11.5316903254, -67.4542168707, 95.5696647599, -29.9496420167};
test_label[4784] = '{-67.4542168707};
test_output[4784] = '{163.023881631};
############ END DEBUG ############*/
test_input[38280:38287] = '{32'h41b6d5b0, 32'h42669a4e, 32'h41d02c90, 32'h41b1e6a9, 32'h4291629f, 32'h423c6afb, 32'h42987a8d, 32'h42940664};
test_label[4785] = '{32'h41b6d5b0};
test_output[4785] = '{32'h42560d73};
/*############ DEBUG ############
test_input[38280:38287] = '{22.8543396747, 57.6506863041, 26.0217593924, 22.2376276177, 72.69261698, 47.1044723694, 76.2393579313, 74.0124778777};
test_label[4785] = '{22.8543396747};
test_output[4785] = '{53.5131324991};
############ END DEBUG ############*/
test_input[38288:38295] = '{32'h411e5322, 32'hc2c76e69, 32'h4289f9a9, 32'hc25e0251, 32'hc2c60059, 32'hc20682ab, 32'hc1d5b240, 32'hc0373a93};
test_label[4786] = '{32'hc20682ab};
test_output[4786] = '{32'h42cd3afe};
/*############ DEBUG ############
test_input[38288:38295] = '{9.89529629225, -99.7156453959, 68.9876169427, -55.5022623842, -99.0006752441, -33.6276039528, -26.7120363947, -2.86295000786};
test_label[4786] = '{-33.6276039528};
test_output[4786] = '{102.615220895};
############ END DEBUG ############*/
test_input[38296:38303] = '{32'hc2a3139a, 32'h426100da, 32'hc1cf6343, 32'hc11a2bb9, 32'hc28f7a5e, 32'h429fe3a9, 32'h429745e2, 32'h42bf99d5};
test_label[4787] = '{32'h42bf99d5};
test_output[4787] = '{32'h340d7475};
/*############ DEBUG ############
test_input[38296:38303] = '{-81.5382854693, 56.250830951, -25.923468396, -9.6356742047, -71.7389958974, 79.9446500712, 75.6364871836, 95.8004529027};
test_label[4787] = '{95.8004529027};
test_output[4787] = '{1.31740151583e-07};
############ END DEBUG ############*/
test_input[38304:38311] = '{32'hc1f55958, 32'h41f43d53, 32'hc22851ce, 32'hc28997a9, 32'hc22427ac, 32'h42aa3974, 32'hc1c24ab6, 32'h4221542c};
test_label[4788] = '{32'hc22851ce};
test_output[4788] = '{32'h42fe625b};
/*############ DEBUG ############
test_input[38304:38311] = '{-30.6686244062, 30.5299437878, -42.0798858152, -68.7962115061, -41.0387411604, 85.112212092, -24.2864795106, 40.332199456};
test_label[4788] = '{-42.0798858152};
test_output[4788] = '{127.192097907};
############ END DEBUG ############*/
test_input[38312:38319] = '{32'hc2a2807f, 32'hc10165f2, 32'hc15bfecb, 32'hc1381238, 32'hc26e2e48, 32'hc2c5c384, 32'h429af689, 32'hc2164e7a};
test_label[4789] = '{32'hc26e2e48};
test_output[4789] = '{32'h430906d6};
/*############ DEBUG ############
test_input[38312:38319] = '{-81.2509690145, -8.08738931344, -13.7497050457, -11.5044478352, -59.5451951633, -98.8818700726, 77.4815144956, -37.5766369996};
test_label[4789] = '{-59.5451951633};
test_output[4789] = '{137.026709659};
############ END DEBUG ############*/
test_input[38320:38327] = '{32'h42ba5647, 32'hc28e4b23, 32'h4230d62d, 32'h427f1cdc, 32'hc28fbc54, 32'h429b3ea8, 32'h40a942a1, 32'h42b78ac8};
test_label[4790] = '{32'h427f1cdc};
test_output[4790] = '{32'h41ece3d6};
/*############ DEBUG ############
test_input[38320:38327] = '{93.1685077773, -71.1467507009, 44.2091548595, 63.7781830205, -71.8678298803, 77.6223770005, 5.28938333568, 91.7710598009};
test_label[4790] = '{63.7781830205};
test_output[4790] = '{29.6112476572};
############ END DEBUG ############*/
test_input[38328:38335] = '{32'h418dc58a, 32'h424c4513, 32'h4221a83a, 32'h41897346, 32'hc2235838, 32'hc1e033e2, 32'hc2b2fdb5, 32'hc2b6866c};
test_label[4791] = '{32'hc1e033e2};
test_output[4791] = '{32'h429e2f85};
/*############ DEBUG ############
test_input[38328:38335] = '{17.721454128, 51.0674566377, 40.4142834273, 17.1812850014, -40.8361525382, -28.0253339567, -89.4955207956, -91.2625434339};
test_label[4791] = '{-28.0253339567};
test_output[4791] = '{79.0928142198};
############ END DEBUG ############*/
test_input[38336:38343] = '{32'hc1cc6de8, 32'hc2a153d9, 32'h42c4a988, 32'h414d523d, 32'hc2bc968e, 32'hc2474fb9, 32'hc2c10057, 32'hc1278021};
test_label[4792] = '{32'hc2bc968e};
test_output[4792] = '{32'h4340a00b};
/*############ DEBUG ############
test_input[38336:38343] = '{-25.5536656372, -80.6637669611, 98.3311127402, 12.8325772776, -94.294053711, -49.8278533799, -96.5006622557, -10.4687812326};
test_label[4792] = '{-94.294053711};
test_output[4792] = '{192.625166451};
############ END DEBUG ############*/
test_input[38344:38351] = '{32'hc08d14b2, 32'h42b0f35c, 32'h424bf96c, 32'hc2b32b9b, 32'hc172b55f, 32'hc11ac363, 32'h3f022785, 32'hc20858cc};
test_label[4793] = '{32'h42b0f35c};
test_output[4793] = '{32'h80000000};
/*############ DEBUG ############
test_input[38344:38351] = '{-4.4087763567, 88.4753136275, 50.9935772667, -89.5851650684, -15.1692798758, -9.672702168, 0.508415549616, -34.0867146539};
test_label[4793] = '{88.4753136275};
test_output[4793] = '{-0.0};
############ END DEBUG ############*/
test_input[38352:38359] = '{32'hc08ec2da, 32'hc20b10a9, 32'hc27b3140, 32'hc2c6853a, 32'hc208a9fb, 32'h428b4f51, 32'h4226ff42, 32'h4185ae49};
test_label[4794] = '{32'hc27b3140};
test_output[4794] = '{32'h430473f8};
/*############ DEBUG ############
test_input[38352:38359] = '{-4.46128556244, -34.7662685613, -62.7980951567, -99.2602083941, -34.1659947787, 69.6549135805, 41.749275295, 16.71010008};
test_label[4794] = '{-62.7980951567};
test_output[4794] = '{132.453008737};
############ END DEBUG ############*/
test_input[38360:38367] = '{32'h406082ff, 32'hc1ff6570, 32'h42790486, 32'hc0cc593d, 32'hc0ed3c05, 32'h428a77ef, 32'h40c6e6fe, 32'hc280d015};
test_label[4795] = '{32'h406082ff};
test_output[4795] = '{32'h42837451};
/*############ DEBUG ############
test_input[38360:38367] = '{3.50799532084, -31.9245297158, 62.2544176377, -6.38589341566, -7.41357641975, 69.2342469196, 6.2156972603, -64.4064084271};
test_label[4795] = '{3.50799532084};
test_output[4795] = '{65.7271816282};
############ END DEBUG ############*/
test_input[38368:38375] = '{32'hc25238dc, 32'hc2689bfe, 32'h41b6b853, 32'hc290beac, 32'h425021a0, 32'hc28dffc5, 32'hc0edaa77, 32'h42653f0d};
test_label[4796] = '{32'hc290beac};
test_output[4796] = '{32'h4301b067};
/*############ DEBUG ############
test_input[38368:38375] = '{-52.5555249437, -58.1523352623, 22.8400019245, -72.3724081195, 52.0328379935, -70.9995531618, -7.42705849201, 57.3115729918};
test_label[4796] = '{-72.3724081195};
test_output[4796] = '{129.689067033};
############ END DEBUG ############*/
test_input[38376:38383] = '{32'h4220ef16, 32'h41d4da98, 32'hc2b0d6af, 32'h42a73d94, 32'hc1f217ad, 32'h40211828, 32'h41da9a4b, 32'hc1d44362};
test_label[4797] = '{32'h4220ef16};
test_output[4797] = '{32'h422d8c12};
/*############ DEBUG ############
test_input[38376:38383] = '{40.2334832232, 26.6067350761, -88.4193022609, 83.620268863, -30.2615605376, 2.51709937608, 27.3253378642, -26.5329025131};
test_label[4797] = '{40.2334832232};
test_output[4797] = '{43.3867856398};
############ END DEBUG ############*/
test_input[38384:38391] = '{32'hc291d834, 32'h3fabf373, 32'h42afea76, 32'h41c8e924, 32'hc15d2e6d, 32'hc299b9b7, 32'h4293c99e, 32'h42905bc8};
test_label[4798] = '{32'hc299b9b7};
test_output[4798] = '{32'h4324d216};
/*############ DEBUG ############
test_input[38384:38391] = '{-72.9222738353, 1.34336700901, 87.9579283902, 25.1138383704, -13.8238342006, -76.8627252448, 73.8937813109, 72.1792614134};
test_label[4798] = '{-76.8627252448};
test_output[4798] = '{164.820654555};
############ END DEBUG ############*/
test_input[38392:38399] = '{32'h42abcc0b, 32'h427376b0, 32'hc1d797f1, 32'h42bb1e73, 32'h42abf876, 32'hc27f6cb7, 32'h41e54bee, 32'h42310939};
test_label[4799] = '{32'h427376b0};
test_output[4799] = '{32'h4202c738};
/*############ DEBUG ############
test_input[38392:38399] = '{85.8985211473, 60.8659051014, -26.9491909656, 93.5594713343, 85.9852777006, -63.8561671324, 28.6620744796, 44.2590078988};
test_label[4799] = '{60.8659051014};
test_output[4799] = '{32.6945501429};
############ END DEBUG ############*/
test_input[38400:38407] = '{32'h42230b5e, 32'hc290ec87, 32'h42858883, 32'hc2ad5e43, 32'hc27be4f2, 32'h429c837d, 32'hc2525736, 32'h42bca864};
test_label[4800] = '{32'h42bca864};
test_output[4800] = '{32'h33e0dd5d};
/*############ DEBUG ############
test_input[38400:38407] = '{40.7610991191, -72.4619668374, 66.7666239435, -86.6841072945, -62.9735793465, 78.2568132526, -52.5851683987, 94.328887173};
test_label[4800] = '{94.328887173};
test_output[4800] = '{1.04710782309e-07};
############ END DEBUG ############*/
test_input[38408:38415] = '{32'h425cc741, 32'hc2360afb, 32'hc1c73298, 32'hc2c5db2b, 32'hc2a62803, 32'h42a06258, 32'hc2bc870d, 32'h426b2082};
test_label[4801] = '{32'hc2360afb};
test_output[4801] = '{32'h42fb67d5};
/*############ DEBUG ############
test_input[38408:38415] = '{55.1945852263, -45.5107225166, -24.8997034882, -98.9280608888, -83.0781461828, 80.1920746869, -94.2637702793, 58.7817478076};
test_label[4801] = '{-45.5107225166};
test_output[4801] = '{125.702797204};
############ END DEBUG ############*/
test_input[38416:38423] = '{32'h3fa7449f, 32'h42930ec8, 32'h41396330, 32'hc0b738ac, 32'hc20ffce5, 32'hc264e9d6, 32'hc157c2f7, 32'hc1c3c2c1};
test_label[4802] = '{32'h41396330};
test_output[4802] = '{32'h4277c4c5};
/*############ DEBUG ############
test_input[38416:38423] = '{1.30678163811, 73.5288721096, 11.5867155326, -5.72566807858, -35.9969660538, -57.2283546005, -13.4850985645, -24.470094639};
test_label[4802] = '{11.5867155326};
test_output[4802] = '{61.942156577};
############ END DEBUG ############*/
test_input[38424:38431] = '{32'hc22568c6, 32'hc2a87038, 32'hc2342f7d, 32'h428aa650, 32'h41956481, 32'hc252cd85, 32'h4170b7dd, 32'h41ce40d7};
test_label[4803] = '{32'hc22568c6};
test_output[4803] = '{32'h42dd5ab2};
/*############ DEBUG ############
test_input[38424:38431] = '{-41.3523164234, -84.2191753768, -45.0463758393, 69.3248260393, 18.6740751095, -52.7007012313, 15.0448888118, 25.7816603612};
test_label[4803] = '{-41.3523164234};
test_output[4803] = '{110.677142463};
############ END DEBUG ############*/
test_input[38432:38439] = '{32'h41d39c29, 32'hc29d0a28, 32'hc2a8dec8, 32'h4148c0eb, 32'hc2a1151e, 32'hc0e4c8e2, 32'hc2741882, 32'hc276e44e};
test_label[4804] = '{32'hc276e44e};
test_output[4804] = '{32'h42b05931};
/*############ DEBUG ############
test_input[38432:38439] = '{26.4512505083, -78.5198394677, -84.4351232861, 12.5470992066, -80.5412413003, -7.14952173873, -61.0239350006, -61.7229533237};
test_label[4804] = '{-61.7229533237};
test_output[4804] = '{88.1742047471};
############ END DEBUG ############*/
test_input[38440:38447] = '{32'hc23b57c3, 32'h3f255c92, 32'hc00a8d14, 32'hc26b2095, 32'hc23264ac, 32'h42b81094, 32'h4285ce43, 32'h4200e396};
test_label[4805] = '{32'hc23264ac};
test_output[4805] = '{32'h4308a175};
/*############ DEBUG ############
test_input[38440:38447] = '{-46.8357066008, 0.64594375551, -2.16486073755, -58.7818183302, -44.5983132396, 92.0323769808, 66.9028563259, 32.2222507124};
test_label[4805] = '{-44.5983132396};
test_output[4805] = '{136.63069022};
############ END DEBUG ############*/
test_input[38448:38455] = '{32'hc1e4f610, 32'h418a3d2e, 32'hc147e56d, 32'h4245061e, 32'hc227f731, 32'h429d85fa, 32'hc298ddfc, 32'h42a859b9};
test_label[4806] = '{32'hc298ddfc};
test_output[4806] = '{32'h43209cfe};
/*############ DEBUG ############
test_input[38448:38455] = '{-28.620148136, 17.2798737971, -12.4935123996, 49.2559750862, -41.9913995306, 78.7616715732, -76.4335603189, 84.1752391579};
test_label[4806] = '{-76.4335603189};
test_output[4806] = '{160.613245295};
############ END DEBUG ############*/
test_input[38456:38463] = '{32'h42bcf3f8, 32'h420b73ae, 32'hc2b98290, 32'h423a0d68, 32'hc2ab9299, 32'hc2c38165, 32'h41840808, 32'h4269445b};
test_label[4807] = '{32'h4269445b};
test_output[4807] = '{32'h4210a394};
/*############ DEBUG ############
test_input[38456:38463] = '{94.4764985419, 34.8629699741, -92.755006906, 46.5130919246, -85.7863220937, -97.75272214, 16.5039221429, 58.3167534185};
test_label[4807] = '{58.3167534185};
test_output[4807] = '{36.1597451234};
############ END DEBUG ############*/
test_input[38464:38471] = '{32'h41b86e9b, 32'hc2536d8b, 32'h428ab15c, 32'hc1efbff0, 32'h422c5179, 32'h41fde32a, 32'hc24aac6b, 32'h424a2ab4};
test_label[4808] = '{32'h424a2ab4};
test_output[4808] = '{32'h41967007};
/*############ DEBUG ############
test_input[38464:38471] = '{23.0540069691, -52.8569766123, 69.3464020834, -29.9687194449, 43.0795636185, 31.7359198816, -50.6683769414, 50.5417007467};
test_label[4808] = '{50.5417007467};
test_output[4808] = '{18.8047013435};
############ END DEBUG ############*/
test_input[38472:38479] = '{32'h41c9e4fe, 32'hc2ab966d, 32'hc19b729d, 32'h3fd846f7, 32'h429448a3, 32'h4270c603, 32'h419bd205, 32'h42ab4969};
test_label[4809] = '{32'hc2ab966d};
test_output[4809] = '{32'h432b6fec};
/*############ DEBUG ############
test_input[38472:38479] = '{25.2368119977, -85.7938039288, -19.4309634659, 1.68966565873, 74.1418669516, 60.1933719522, 19.4775493447, 85.6433788778};
test_label[4809] = '{-85.7938039288};
test_output[4809] = '{171.437192921};
############ END DEBUG ############*/
test_input[38480:38487] = '{32'hc19aa15f, 32'h428ff3c9, 32'h41b7b54c, 32'hc24cc4be, 32'h4245f5f4, 32'h428cde91, 32'hc1caf779, 32'hc209f723};
test_label[4810] = '{32'hc24cc4be};
test_output[4810] = '{32'h42f6b979};
/*############ DEBUG ############
test_input[38480:38487] = '{-19.3287941442, 71.9761447375, 22.9635232153, -51.1921300077, 49.4901884875, 70.4347003981, -25.3708363587, -34.4913462991};
test_label[4810] = '{-51.1921300077};
test_output[4810] = '{123.362254486};
############ END DEBUG ############*/
test_input[38488:38495] = '{32'hc20887ea, 32'h40fbfacb, 32'h41aa0b67, 32'hc220e750, 32'hc25f4ea1, 32'h4147007f, 32'h42c33fdb, 32'hc28da01c};
test_label[4811] = '{32'h40fbfacb};
test_output[4811] = '{32'h42b3802e};
/*############ DEBUG ############
test_input[38488:38495] = '{-34.1327274213, 7.87436422665, 21.2555680298, -40.2258897223, -55.8267844707, 12.4376214728, 97.6247150734, -70.8127134425};
test_label[4811] = '{7.87436422665};
test_output[4811] = '{89.7503508467};
############ END DEBUG ############*/
test_input[38496:38503] = '{32'h429b85c7, 32'h41a16ecd, 32'h4273ff09, 32'hc2144d58, 32'hc2646e0c, 32'hc0eae0ef, 32'hc14a15c0, 32'h4290b453};
test_label[4812] = '{32'hc2646e0c};
test_output[4812] = '{32'h4306df8b};
/*############ DEBUG ############
test_input[38496:38503] = '{77.7612818089, 20.1791014693, 60.9990576473, -37.0755301706, -57.1074675797, -7.33995776961, -12.6303098017, 72.3521982903};
test_label[4812] = '{-57.1074675797};
test_output[4812] = '{134.873215195};
############ END DEBUG ############*/
test_input[38504:38511] = '{32'hc2952910, 32'hc245b0bb, 32'h405590cc, 32'h4243b969, 32'h4060b1fd, 32'hc0fb1ba7, 32'h42964d24, 32'hc2acf2d7};
test_label[4813] = '{32'hc2952910};
test_output[4813] = '{32'h4315bb1a};
/*############ DEBUG ############
test_input[38504:38511] = '{-74.5801995938, -49.422589307, 3.33696276119, 48.9310650971, 3.5108634412, -7.84712561535, 75.1506671791, -86.4742934825};
test_label[4813] = '{-74.5801995938};
test_output[4813] = '{149.730866773};
############ END DEBUG ############*/
test_input[38512:38519] = '{32'h4144b9a2, 32'hc273f064, 32'hc2a865a8, 32'hc26377cd, 32'hc2333f59, 32'h420c5e31, 32'hc2a95cde, 32'h41df769b};
test_label[4814] = '{32'hc2333f59};
test_output[4814] = '{32'h429fcf2b};
/*############ DEBUG ############
test_input[38512:38519] = '{12.2953208937, -60.9847583673, -84.1985474833, -56.8669933066, -44.8118644863, 35.0919833489, -84.6813806066, 27.9329129361};
test_label[4814] = '{-44.8118644863};
test_output[4814] = '{79.9046253103};
############ END DEBUG ############*/
test_input[38520:38527] = '{32'h42bec23a, 32'h42046658, 32'h42678262, 32'hc232141e, 32'hc2897492, 32'hc2c5310b, 32'hc1e4803d, 32'h42435374};
test_label[4815] = '{32'hc1e4803d};
test_output[4815] = '{32'h42f7e249};
/*############ DEBUG ############
test_input[38520:38527] = '{95.379346876, 33.0999435743, 57.8773265526, -44.5196463386, -68.7276741207, -98.5957889337, -28.5626154124, 48.8314960846};
test_label[4815] = '{-28.5626154124};
test_output[4815] = '{123.941962288};
############ END DEBUG ############*/
test_input[38528:38535] = '{32'h424482ca, 32'hc21634f9, 32'h42bdca3c, 32'hc0836e2a, 32'hc270abdd, 32'hc2118d4e, 32'hc2b299ae, 32'h421afa4a};
test_label[4816] = '{32'hc270abdd};
test_output[4816] = '{32'h431b1015};
/*############ DEBUG ############
test_input[38528:38535] = '{49.1277240446, -37.5517306758, 94.8949908903, -4.10719764433, -60.167834405, -36.3879938956, -89.3001548516, 38.7444212041};
test_label[4816] = '{-60.167834405};
test_output[4816] = '{155.062825295};
############ END DEBUG ############*/
test_input[38536:38543] = '{32'hc206d869, 32'h41be82a6, 32'h429313b2, 32'hc2aa43ac, 32'h428ea2b8, 32'h42665395, 32'hc204d2da, 32'h4223fa93};
test_label[4817] = '{32'hc204d2da};
test_output[4817] = '{32'h42d5b1e1};
/*############ DEBUG ############
test_input[38536:38543] = '{-33.7113395668, 23.813793054, 73.5384677458, -85.1321695086, 71.3178127789, 57.581624741, -33.2059088489, 40.9947013079};
test_label[4817] = '{-33.2059088489};
test_output[4817] = '{106.847418728};
############ END DEBUG ############*/
test_input[38544:38551] = '{32'h42bef9a9, 32'hc26bc465, 32'h40cda75c, 32'h42864412, 32'h42908bf7, 32'hc188ad83, 32'hc28cc049, 32'hc16260c7};
test_label[4818] = '{32'h42bef9a9};
test_output[4818] = '{32'h2eb73540};
/*############ DEBUG ############
test_input[38544:38551] = '{95.4876208819, -58.9417918055, 6.42667937791, 67.1329488393, 72.2733700787, -17.0847216896, -70.375555157, -14.148627039};
test_label[4818] = '{95.4876208819};
test_output[4818] = '{8.33133562174e-11};
############ END DEBUG ############*/
test_input[38552:38559] = '{32'hc2abd4b3, 32'hc298a2bb, 32'h4280e8dc, 32'hc2b311e2, 32'hc29d5b7c, 32'h423fe147, 32'h4184b8fc, 32'h4200534b};
test_label[4819] = '{32'hc2b311e2};
test_output[4819] = '{32'h4319fd5f};
/*############ DEBUG ############
test_input[38552:38559] = '{-85.9154281524, -76.3178365466, 64.4548011191, -89.5349306611, -78.6786780588, 47.9699992897, 16.5903250056, 32.0813390816};
test_label[4819] = '{-89.5349306611};
test_output[4819] = '{153.98973185};
############ END DEBUG ############*/
test_input[38560:38567] = '{32'hc21cb3b7, 32'h42c4b5bd, 32'h42078bbf, 32'h419015ba, 32'h403f5c0b, 32'h41bc968f, 32'hc211aedb, 32'h428ce65f};
test_label[4820] = '{32'h42c4b5bd};
test_output[4820] = '{32'h2b560000};
/*############ DEBUG ############
test_input[38560:38567] = '{-39.1755042691, 98.3549583713, 33.8864694497, 18.0106082217, 2.98999293295, 23.5735156497, -36.420758609, 70.4499449629};
test_label[4820] = '{98.3549583713};
test_output[4820] = '{7.60280727264e-13};
############ END DEBUG ############*/
test_input[38568:38575] = '{32'hc209bd26, 32'hc24fa379, 32'h42955ca2, 32'h41705004, 32'hc1b27fff, 32'h42aca8fe, 32'hc1af0690, 32'h424974a5};
test_label[4821] = '{32'h41705004};
test_output[4821] = '{32'h428e9efe};
/*############ DEBUG ############
test_input[38568:38575] = '{-34.4347143504, -51.909642358, 74.6809218535, 15.0195352812, -22.3124989929, 86.3300615168, -21.8782045099, 50.3639120985};
test_label[4821] = '{15.0195352812};
test_output[4821] = '{71.3105349621};
############ END DEBUG ############*/
test_input[38576:38583] = '{32'hc1ee7d92, 32'h428494d8, 32'h4282be43, 32'hc217e869, 32'hc2241234, 32'hc2ba3519, 32'h42ae2b54, 32'hc2bd67a9};
test_label[4822] = '{32'h428494d8};
test_output[4822] = '{32'h41a659f0};
/*############ DEBUG ############
test_input[38576:38583] = '{-29.8113140322, 66.290706636, 65.3716064861, -37.9769624122, -41.0177754585, -93.103707428, 87.0846217701, -94.7024603773};
test_label[4822] = '{66.290706636};
test_output[4822] = '{20.7939151353};
############ END DEBUG ############*/
test_input[38584:38591] = '{32'h42b8cc2d, 32'h426b280f, 32'h429013cb, 32'h41fe57d6, 32'hc2213f6c, 32'hc2847c74, 32'h42ab9d06, 32'h428cb52f};
test_label[4823] = '{32'h42b8cc2d};
test_output[4823] = '{32'h3ab39951};
/*############ DEBUG ############
test_input[38584:38591] = '{92.3987773512, 58.7891205665, 72.0386558447, 31.7928893446, -40.3119350384, -66.2430759546, 85.8066852194, 70.3538732181};
test_label[4823] = '{92.3987773512};
test_output[4823] = '{0.00137023080541};
############ END DEBUG ############*/
test_input[38592:38599] = '{32'hc26fd7d7, 32'h4260d122, 32'hc104dd06, 32'hc219dc05, 32'h4097e57e, 32'hc1b39bcc, 32'h42ac8ecf, 32'hc1b75111};
test_label[4824] = '{32'h4260d122};
test_output[4824] = '{32'h41f098fa};
/*############ DEBUG ############
test_input[38592:38599] = '{-59.9607802915, 56.204229621, -8.30396040297, -38.4648640813, 4.74676440409, -22.4510717981, 86.2789248422, -22.9145827331};
test_label[4824] = '{56.204229621};
test_output[4824] = '{30.0746952212};
############ END DEBUG ############*/
test_input[38600:38607] = '{32'h42c0d09b, 32'h428775ef, 32'hc25d9975, 32'hc28a7be2, 32'hc1853d13, 32'h42bbaf54, 32'h42679a8d, 32'h3dd23a4d};
test_label[4825] = '{32'hc1853d13};
test_output[4825] = '{32'h42e245d0};
/*############ DEBUG ############
test_input[38600:38607] = '{96.4074291655, 67.7303407464, -55.3998621151, -69.2419607764, -16.6548210601, 93.842436921, 57.9009276242, 0.102650261213};
test_label[4825] = '{-16.6548210601};
test_output[4825] = '{113.136355134};
############ END DEBUG ############*/
test_input[38608:38615] = '{32'hc130dd07, 32'hc20b2a24, 32'h41939f17, 32'h41b559c4, 32'h4277c634, 32'h40a11930, 32'hc262478f, 32'h4295b838};
test_label[4826] = '{32'hc20b2a24};
test_output[4826] = '{32'h42db4d4a};
/*############ DEBUG ############
test_input[38608:38615] = '{-11.0539614925, -34.7911545891, 18.4526806513, 22.668831525, 61.9435572547, 5.03432465871, -56.5698795329, 74.8597989806};
test_label[4826] = '{-34.7911545891};
test_output[4826] = '{109.650956028};
############ END DEBUG ############*/
test_input[38616:38623] = '{32'h41f12586, 32'hc2bd5182, 32'hc24d5013, 32'hc1dbb7fc, 32'h4118f973, 32'h42ad688a, 32'h42822e6f, 32'h427f7815};
test_label[4827] = '{32'h4118f973};
test_output[4827] = '{32'h429a495c};
/*############ DEBUG ############
test_input[38616:38623] = '{30.1433226137, -94.659193701, -51.3281978095, -27.4648354586, 9.56090107672, 86.7041811423, 65.0906913882, 63.8672685056};
test_label[4827] = '{9.56090107672};
test_output[4827] = '{77.1432800661};
############ END DEBUG ############*/
test_input[38624:38631] = '{32'h41888978, 32'hbfe025e3, 32'hc1ad82d9, 32'hc2afc16a, 32'h415adcce, 32'hc206c4d8, 32'h428e7a9a, 32'hc16c339f};
test_label[4828] = '{32'hbfe025e3};
test_output[4828] = '{32'h4291fb31};
/*############ DEBUG ############
test_input[38624:38631] = '{17.0671236793, -1.75115622892, -21.6888906762, -87.8777643468, 13.6789070662, -33.6922287949, 71.2394534326, -14.7626028814};
test_label[4828] = '{-1.75115622892};
test_output[4828] = '{72.9906096615};
############ END DEBUG ############*/
test_input[38632:38639] = '{32'hc246c56f, 32'h42721f5c, 32'h429a0ad6, 32'h42660fa9, 32'hc2c13337, 32'hc2ada31d, 32'hc1036951, 32'h426ef247};
test_label[4829] = '{32'h42660fa9};
test_output[4829] = '{32'h419c0c07};
/*############ DEBUG ############
test_input[38632:38639] = '{-49.692806008, 60.530625881, 77.0211655741, 57.5152928903, -96.6000254943, -86.8185800808, -8.21321187571, 59.7365978607};
test_label[4829] = '{57.5152928903};
test_output[4829] = '{19.5058727872};
############ END DEBUG ############*/
test_input[38640:38647] = '{32'hc20b7089, 32'hc2ad015d, 32'hc22cb50c, 32'h3f5e0169, 32'hc247b972, 32'h42384e1a, 32'h406b5342, 32'h42003a9e};
test_label[4830] = '{32'h42384e1a};
test_output[4830] = '{32'h355b0130};
/*############ DEBUG ############
test_input[38640:38647] = '{-34.8598962402, -86.502659496, -43.1768046653, 0.86720902091, -49.931097335, 46.0762724451, 3.6769566564, 32.0572447064};
test_label[4830] = '{46.0762724451};
test_output[4830] = '{8.15855854285e-07};
############ END DEBUG ############*/
test_input[38648:38655] = '{32'hc278a5c2, 32'hc1a2e297, 32'h42c4f61b, 32'hc1fe2fa2, 32'hc1fac5fb, 32'h42be50ea, 32'h40e0b71b, 32'h414c1ac5};
test_label[4831] = '{32'h42be50ea};
test_output[4831] = '{32'h4056ea7e};
/*############ DEBUG ############
test_input[38648:38655] = '{-62.1618714308, -20.360639991, 98.4806729056, -31.7732589529, -31.3466700747, 95.1580332143, 7.02235165591, 12.7565356551};
test_label[4831] = '{95.1580332143};
test_output[4831] = '{3.35806235996};
############ END DEBUG ############*/
test_input[38656:38663] = '{32'h429d74ae, 32'h41e78562, 32'hbfc2121d, 32'hc158019c, 32'h42830e0c, 32'hc24f8330, 32'h425b5f21, 32'hc280142b};
test_label[4832] = '{32'h429d74ae};
test_output[4832] = '{32'h35f846c4};
/*############ DEBUG ############
test_input[38656:38663] = '{78.727888005, 28.940127827, -1.5161777912, -13.5003924918, 65.527434892, -51.878112481, 54.8428974433, -64.0393928823};
test_label[4832] = '{78.727888005};
test_output[4832] = '{1.84980349785e-06};
############ END DEBUG ############*/
test_input[38664:38671] = '{32'h42c79e02, 32'h4046a54d, 32'h42a06c8c, 32'h42979789, 32'hc233b7be, 32'hc291c5b6, 32'hc23af4cc, 32'h42b92bab};
test_label[4833] = '{32'h42979789};
test_output[4833] = '{32'h41c01b63};
/*############ DEBUG ############
test_input[38664:38671] = '{99.8086084483, 3.10383917927, 80.2120069466, 75.7959659127, -44.9294366838, -72.8861511206, -46.7390590759, 92.585287104};
test_label[4833] = '{75.7959659127};
test_output[4833] = '{24.0133716487};
############ END DEBUG ############*/
test_input[38672:38679] = '{32'h421c9b07, 32'hc09df28b, 32'h42b2ba7f, 32'hc2c7ecf3, 32'hc0cff13c, 32'h41f6a003, 32'h427a38d3, 32'hc14c61b9};
test_label[4834] = '{32'hc14c61b9};
test_output[4834] = '{32'h42cc46b6};
/*############ DEBUG ############
test_input[38672:38679] = '{39.1513940109, -4.93585710219, 89.3642501253, -99.9627882841, -6.49819766926, 30.8281307604, 62.55549312, -12.7738582469};
test_label[4834] = '{-12.7738582469};
test_output[4834] = '{102.138108372};
############ END DEBUG ############*/
test_input[38680:38687] = '{32'hc270755e, 32'h421e9aa1, 32'h42b29482, 32'h424bc9ee, 32'h41f5cbc2, 32'hc1297108, 32'h4184ac27, 32'h42469fbe};
test_label[4835] = '{32'h4184ac27};
test_output[4835] = '{32'h42916978};
/*############ DEBUG ############
test_input[38680:38687] = '{-60.1146150579, 39.6510058733, 89.2900545287, 50.9471959213, 30.7244902081, -10.5900957646, 16.5840593668, 49.65599859};
test_label[4835] = '{16.5840593668};
test_output[4835] = '{72.7059951619};
############ END DEBUG ############*/
test_input[38688:38695] = '{32'h42a4ec6f, 32'h428bea71, 32'h42aa69b2, 32'hc22457c7, 32'h41f3ca1a, 32'h42bd485d, 32'h428985f3, 32'hc2ada57c};
test_label[4836] = '{32'h42aa69b2};
test_output[4836] = '{32'h4116f5b0};
/*############ DEBUG ############
test_input[38688:38695] = '{82.4617850751, 69.9578969987, 85.2064384314, -41.0857204294, 30.4736823192, 94.6413356524, 68.7616209385, -86.823215346};
test_label[4836] = '{85.2064384314};
test_output[4836] = '{9.43498223881};
############ END DEBUG ############*/
test_input[38696:38703] = '{32'hc211f340, 32'hc213aebb, 32'hc28f0ede, 32'h419758e6, 32'hc20efa69, 32'hc1899554, 32'h4136b919, 32'hc2695c00};
test_label[4837] = '{32'hc28f0ede};
test_output[4837] = '{32'h42b4e560};
/*############ DEBUG ############
test_input[38696:38703] = '{-36.4875496447, -36.9206338079, -71.5290347253, 18.918407858, -35.744539717, -17.1979148404, 11.4201901869, -58.3398433767};
test_label[4837] = '{-71.5290347253};
test_output[4837] = '{90.4479965009};
############ END DEBUG ############*/
test_input[38704:38711] = '{32'h42a32799, 32'hc20d7ab4, 32'hc27dffda, 32'hc1ce8ba0, 32'hc20a619d, 32'h40e3340d, 32'hc18ef33b, 32'h414269c3};
test_label[4838] = '{32'h414269c3};
test_output[4838] = '{32'h428ada61};
/*############ DEBUG ############
test_input[38704:38711] = '{81.5773400798, -35.3698265685, -63.4998549766, -25.8181760832, -34.5953243007, 7.10010387549, -17.8687641538, 12.1508204839};
test_label[4838] = '{12.1508204839};
test_output[4838] = '{69.4265195959};
############ END DEBUG ############*/
test_input[38712:38719] = '{32'h411841da, 32'h42c4eb74, 32'hc1698730, 32'hc2bdb1da, 32'hc2a02981, 32'h423f6ffb, 32'h41d397b2, 32'h42283325};
test_label[4839] = '{32'h42283325};
test_output[4839] = '{32'h4261a3c4};
/*############ DEBUG ############
test_input[38712:38719] = '{9.51607668465, 98.4598730119, -14.595504672, -94.8473676868, -80.0810616415, 47.8593560229, 26.449070214, 42.0499471356};
test_label[4839] = '{42.0499471356};
test_output[4839] = '{56.4099258762};
############ END DEBUG ############*/
test_input[38720:38727] = '{32'hc1b4cd94, 32'hc108d9b7, 32'h4210ef16, 32'h41c67871, 32'h4154bfcb, 32'h41afb525, 32'hc28743d4, 32'hc2c5235b};
test_label[4840] = '{32'h4210ef16};
test_output[4840] = '{32'h3741e6e6};
/*############ DEBUG ############
test_input[38720:38727] = '{-22.6003802689, -8.55315350435, 36.2334808234, 24.8088100173, 13.2968242263, 21.9634491536, -67.6324734614, -98.5690522864};
test_label[4840] = '{36.2334808234};
test_output[4840] = '{1.15574568319e-05};
############ END DEBUG ############*/
test_input[38728:38735] = '{32'hbf2a8d9f, 32'hc254de74, 32'hc29e188b, 32'h422e83c7, 32'h4297449d, 32'h40a77254, 32'hc0fc4da2, 32'h4031a487};
test_label[4841] = '{32'h4031a487};
test_output[4841] = '{32'h4291b778};
/*############ DEBUG ############
test_input[38728:38735] = '{-0.666223486686, -53.2172397022, -79.0479321381, 43.6286898091, 75.6340077436, 5.23270629149, -7.8844766626, 2.77566686246};
test_label[4841] = '{2.77566686246};
test_output[4841] = '{72.8583408811};
############ END DEBUG ############*/
test_input[38736:38743] = '{32'hc272bce4, 32'h429a044a, 32'hc247750e, 32'h4220f0f8, 32'hc2838ad1, 32'hc0901ee1, 32'hc297fea4, 32'hc18040df};
test_label[4842] = '{32'hc272bce4};
test_output[4842] = '{32'h4309b15e};
/*############ DEBUG ############
test_input[38736:38743] = '{-60.684463625, 77.0083766067, -49.8643115691, 40.2353215067, -65.7711261108, -4.5037693338, -75.9973430232, -16.0316751294};
test_label[4842] = '{-60.684463625};
test_output[4842] = '{137.692840232};
############ END DEBUG ############*/
test_input[38744:38751] = '{32'hc1de478b, 32'hc2516fc0, 32'h4233bc2a, 32'hc2c02428, 32'hc1fa4e21, 32'h41a78114, 32'hc1b12269, 32'h41d4fe58};
test_label[4843] = '{32'hc1de478b};
test_output[4843] = '{32'h42916ff8};
/*############ DEBUG ############
test_input[38744:38751] = '{-27.7849329557, -52.3591303801, 44.9337522483, -96.0706187933, -31.2881493993, 20.9380271323, -22.1418026946, 26.6241910758};
test_label[4843] = '{-27.7849329557};
test_output[4843] = '{72.7186852152};
############ END DEBUG ############*/
test_input[38752:38759] = '{32'hc11929da, 32'hc25e1829, 32'h426b71a3, 32'hc21879ca, 32'hc2a85d4b, 32'h427fcc8b, 32'hc2556d65, 32'hc263404a};
test_label[4844] = '{32'hc11929da};
test_output[4844] = '{32'h42930ea6};
/*############ DEBUG ############
test_input[38752:38759] = '{-9.57271733916, -55.5235933705, 58.8609729347, -38.1189332742, -84.1822126598, 63.9497489984, -53.35682959, -56.8127812908};
test_label[4844] = '{-9.57271733916};
test_output[4844] = '{73.5286129697};
############ END DEBUG ############*/
test_input[38760:38767] = '{32'h42917267, 32'hc1af67bf, 32'hc2c1313a, 32'hc280e5b0, 32'hc2ad75b5, 32'hc2055010, 32'hc1e92b4c, 32'hc221a814};
test_label[4845] = '{32'hc2055010};
test_output[4845] = '{32'h42d41a6f};
/*############ DEBUG ############
test_input[38760:38767] = '{72.7234438312, -21.925656975, -96.5961460529, -64.4486114353, -86.7298948784, -33.3281861837, -29.1461416845, -40.4141372408};
test_label[4845] = '{-33.3281861837};
test_output[4845] = '{106.051630015};
############ END DEBUG ############*/
test_input[38768:38775] = '{32'h413d1a03, 32'hc2b03698, 32'h429b186b, 32'h42a088ba, 32'h42bc782c, 32'hc1dabe83, 32'hc2b48354, 32'hc29f060a};
test_label[4846] = '{32'h429b186b};
test_output[4846] = '{32'h41857f02};
/*############ DEBUG ############
test_input[38768:38775] = '{11.8188503702, -88.1066291426, 77.5476924523, 80.2670402998, 94.2347075819, -27.3430242358, -90.2564983205, -79.5117974376};
test_label[4846] = '{77.5476924523};
test_output[4846] = '{16.687016045};
############ END DEBUG ############*/
test_input[38776:38783] = '{32'h421ae197, 32'hc22285f5, 32'hc2c7824b, 32'h42409347, 32'hc2c465a5, 32'hc21d8e52, 32'h4289bb19, 32'hc2900242};
test_label[4847] = '{32'h421ae197};
test_output[4847] = '{32'h41f12936};
/*############ DEBUG ############
test_input[38776:38783] = '{38.7203014441, -40.6308179851, -99.7544803305, 48.1438262872, -98.1985236947, -39.3889855249, 68.8654242449, -72.0044101667};
test_label[4847] = '{38.7203014441};
test_output[4847] = '{30.1451228017};
############ END DEBUG ############*/
test_input[38784:38791] = '{32'hc22d13a3, 32'hc1dea4d0, 32'h41a28da4, 32'hc2830acd, 32'hbf2e383e, 32'hc213ac95, 32'hc2a06d27, 32'hc2c70491};
test_label[4848] = '{32'hbf2e383e};
test_output[4848] = '{32'h41a7ff66};
/*############ DEBUG ############
test_input[38784:38791] = '{-43.2691773706, -27.8304747239, 20.3191607766, -65.5210957759, -0.680545695607, -36.9185360697, -80.21319163, -99.5089210006};
test_label[4848] = '{-0.680545695607};
test_output[4848] = '{20.9997064729};
############ END DEBUG ############*/
test_input[38792:38799] = '{32'hc0bd84c7, 32'hc16a3b25, 32'h4292b72b, 32'hc26092fe, 32'hc25ab29f, 32'hc2a13bdf, 32'hc29f8b3c, 32'hc021ba15};
test_label[4849] = '{32'hc2a13bdf};
test_output[4849] = '{32'h4319f985};
/*############ DEBUG ############
test_input[38792:38799] = '{-5.92245812003, -14.6394391115, 73.3577515221, -56.143548563, -54.6744331397, -80.6169325459, -79.7719452351, -2.5269825552};
test_label[4849] = '{-80.6169325459};
test_output[4849] = '{153.974684068};
############ END DEBUG ############*/
test_input[38800:38807] = '{32'h42b22db3, 32'h41f5e3d9, 32'hc1d07183, 32'hc1c0d023, 32'hc22ab79d, 32'hc13a649f, 32'hc1a4e2a1, 32'h4103cffb};
test_label[4850] = '{32'h41f5e3d9};
test_output[4850] = '{32'h42696979};
/*############ DEBUG ############
test_input[38800:38807] = '{89.0892530514, 30.7362538972, -26.0554258825, -24.1016294325, -42.6793081747, -11.6495653534, -20.6106579774, 8.23827676052};
test_label[4850] = '{30.7362538972};
test_output[4850] = '{58.3529991542};
############ END DEBUG ############*/
test_input[38808:38815] = '{32'h42877ff2, 32'h42bdef57, 32'h426d1a7d, 32'h42999f9b, 32'hc20c7225, 32'hc1a30fda, 32'hc2a4e46f, 32'hc267329a};
test_label[4851] = '{32'hc267329a};
test_output[4851] = '{32'h4318c452};
/*############ DEBUG ############
test_input[38808:38815] = '{67.74989566, 94.9674629928, 59.2758684191, 76.8117321439, -35.1114696159, -20.3827393889, -82.4461576872, -57.7994142986};
test_label[4851] = '{-57.7994142986};
test_output[4851] = '{152.766877304};
############ END DEBUG ############*/
test_input[38816:38823] = '{32'h4208b5fd, 32'hc234824d, 32'hc2562f6f, 32'hc1ff7a41, 32'hc2c477d3, 32'hc2bfc1ba, 32'hc216c642, 32'hc23ea178};
test_label[4852] = '{32'hc2bfc1ba};
test_output[4852] = '{32'h43020e5c};
/*############ DEBUG ############
test_input[38816:38823] = '{34.1777229476, -45.1272452964, -53.546320082, -31.9346936676, -98.2340283038, -95.878369912, -37.6936098686, -47.6576831613};
test_label[4852] = '{-95.878369912};
test_output[4852] = '{130.05609286};
############ END DEBUG ############*/
test_input[38824:38831] = '{32'h42869d9c, 32'h41f9e0f5, 32'hbf92a75a, 32'h42c16b57, 32'h410a226d, 32'hc283f716, 32'h4288e780, 32'hc25e308b};
test_label[4853] = '{32'hc25e308b};
test_output[4853] = '{32'h431841ce};
/*############ DEBUG ############
test_input[38824:38831] = '{67.3078304009, 31.2348413836, -1.14573219943, 96.70964651, 8.63340514347, -65.9825874506, 68.4521460322, -55.547403504};
test_label[4853] = '{-55.547403504};
test_output[4853] = '{152.257050014};
############ END DEBUG ############*/
test_input[38832:38839] = '{32'h42b3478f, 32'h41cf0303, 32'hc19150df, 32'h41b25585, 32'hc0edb369, 32'h4206fdd8, 32'h424714df, 32'h41b3f6e6};
test_label[4854] = '{32'h424714df};
test_output[4854] = '{32'h421f7a3f};
/*############ DEBUG ############
test_input[38832:38839] = '{89.6397650774, 25.8764707895, -18.1644875753, 22.2917572921, -7.42815041685, 33.7478954705, 49.7703831454, 22.4955557714};
test_label[4854] = '{49.7703831454};
test_output[4854] = '{39.869381932};
############ END DEBUG ############*/
test_input[38840:38847] = '{32'hc295b0b2, 32'h4110c88d, 32'hc2a0e02e, 32'hc1d26c9a, 32'h41a01b78, 32'h40fa49ef, 32'hc0bbf612, 32'hc2b151b4};
test_label[4855] = '{32'hc2b151b4};
test_output[4855] = '{32'h42d95895};
/*############ DEBUG ############
test_input[38840:38847] = '{-74.8451043719, 9.04896218126, -80.4378494445, -26.3030275958, 20.013412335, 7.82152513255, -5.87378767538, -88.6595732856};
test_label[4855] = '{-88.6595732856};
test_output[4855] = '{108.673007998};
############ END DEBUG ############*/
test_input[38848:38855] = '{32'hc2142db2, 32'hc2a79bcb, 32'hc211d60e, 32'hc2b432d4, 32'h422b2874, 32'hc2216d0c, 32'hc2ac6dee, 32'hc255315e};
test_label[4856] = '{32'hc2a79bcb};
test_output[4856] = '{32'h42fd3005};
/*############ DEBUG ############
test_input[38848:38855] = '{-37.044624572, -83.8042853413, -36.4590394345, -90.0992710358, 42.7895053449, -40.3564903518, -86.2147070166, -53.2982117862};
test_label[4856] = '{-83.8042853413};
test_output[4856] = '{126.593790686};
############ END DEBUG ############*/
test_input[38856:38863] = '{32'h40496b0b, 32'h412ce8dd, 32'hc297b942, 32'hc2993091, 32'hbf588018, 32'h4229a764, 32'hc24efbc6, 32'h4230b52b};
test_label[4857] = '{32'h4230b52b};
test_output[4857] = '{32'h3e220a9b};
/*############ DEBUG ############
test_input[38856:38863] = '{3.14715832525, 10.8068511989, -75.8618313211, -76.5948592604, -0.84570457912, 42.4134684738, -51.7458716433, 44.1769233399};
test_label[4857] = '{44.1769233399};
test_output[4857] = '{0.158243576011};
############ END DEBUG ############*/
test_input[38864:38871] = '{32'h426e6be2, 32'h42c32ea9, 32'hc2a9b77f, 32'hc1dfae62, 32'hc2199bf2, 32'h429139fb, 32'h40902e1b, 32'h41c9715f};
test_label[4858] = '{32'hc2199bf2};
test_output[4858] = '{32'h4307fe51};
/*############ DEBUG ############
test_input[38864:38871] = '{59.6053560432, 97.5911332799, -84.8583873395, -27.9601483182, -38.4022916665, 72.6132425321, 4.50562787072, 25.1803575801};
test_label[4858] = '{-38.4022916665};
test_output[4858] = '{135.993424946};
############ END DEBUG ############*/
test_input[38872:38879] = '{32'h412a4760, 32'hc29b6972, 32'h403eb1ae, 32'h4222f45b, 32'h412bd173, 32'hc18e6d69, 32'h42bab97f, 32'hc06380a8};
test_label[4859] = '{32'h403eb1ae};
test_output[4859] = '{32'h42b4c3f1};
/*############ DEBUG ############
test_input[38872:38879] = '{10.6424254746, -77.7059472589, 2.97959463553, 40.7386292199, 10.7386354884, -17.8034224179, 93.3622932652, -3.55472746712};
test_label[4859] = '{2.97959463553};
test_output[4859] = '{90.3826986297};
############ END DEBUG ############*/
test_input[38880:38887] = '{32'hc2057a41, 32'hc298983c, 32'hc191392e, 32'hc222e159, 32'hc2065c9d, 32'h4242091d, 32'h42aa2ca0, 32'h41323f37};
test_label[4860] = '{32'h4242091d};
test_output[4860] = '{32'h42125023};
/*############ DEBUG ############
test_input[38880:38887] = '{-33.3693893147, -76.2973345395, -18.1529191785, -40.720065208, -33.5904413811, 48.5088992957, 85.0871588855, 11.1404337018};
test_label[4860] = '{48.5088992957};
test_output[4860] = '{36.5782595898};
############ END DEBUG ############*/
test_input[38888:38895] = '{32'h42c3c573, 32'h41ffb7ff, 32'h40f56c8d, 32'h417174b9, 32'h425610fd, 32'h4131ba01, 32'hc2ab5e61, 32'hc290e1e6};
test_label[4861] = '{32'h41ffb7ff};
test_output[4861] = '{32'h4283d774};
/*############ DEBUG ############
test_input[38888:38895] = '{97.8856460058, 31.9648422669, 7.66950059479, 15.0909968873, 53.5165907498, 11.1079115539, -85.6843354141, -72.4412102478};
test_label[4861] = '{31.9648422669};
test_output[4861] = '{65.9208037389};
############ END DEBUG ############*/
test_input[38896:38903] = '{32'hc2828aa5, 32'h40149d79, 32'h42a91420, 32'h41d01792, 32'h421a3031, 32'hc24da484, 32'hc1fdc2e8, 32'hc0abe46b};
test_label[4862] = '{32'hc24da484};
test_output[4862] = '{32'h4307f331};
/*############ DEBUG ############
test_input[38896:38903] = '{-65.2707915592, 2.32211148637, 84.5393058469, 26.0115097188, 38.5470615766, -51.4106607693, -31.7201699944, -5.37163297588};
test_label[4862] = '{-51.4106607693};
test_output[4862] = '{135.949966616};
############ END DEBUG ############*/
test_input[38904:38911] = '{32'h429da0f1, 32'h426fc1a6, 32'h42abdce2, 32'hc2b6cc91, 32'h422dc246, 32'hc212d42d, 32'hc289d536, 32'h41de7110};
test_label[4863] = '{32'h422dc246};
test_output[4863] = '{32'h4229f852};
/*############ DEBUG ############
test_input[38904:38911] = '{78.8143360088, 59.9391115307, 85.9314089493, -91.3995473331, 43.439719851, -36.7072027789, -68.9164261824, 27.8052055824};
test_label[4863] = '{43.439719851};
test_output[4863] = '{42.4924999071};
############ END DEBUG ############*/
test_input[38912:38919] = '{32'h429de69b, 32'h42b82d74, 32'h428c62f8, 32'hc066a912, 32'hc2a1ea0c, 32'h42841d28, 32'h42a8ea69, 32'h42b8c8da};
test_label[4864] = '{32'h428c62f8};
test_output[4864] = '{32'h41b60437};
/*############ DEBUG ############
test_input[38912:38919] = '{78.9504024429, 92.0887736353, 70.1932983451, -3.60406923703, -80.9571255585, 66.0569431791, 84.4578313159, 92.3922886484};
test_label[4864] = '{70.1932983451};
test_output[4864] = '{22.7520580973};
############ END DEBUG ############*/
test_input[38920:38927] = '{32'hc2b63abd, 32'hc2676fd2, 32'h41b0a30b, 32'h42ac9c07, 32'h4089e4c2, 32'h3f5ca2e2, 32'h41a43815, 32'hc240c8d3};
test_label[4865] = '{32'h41a43815};
test_output[4865] = '{32'h42838e02};
/*############ DEBUG ############
test_input[38920:38927] = '{-91.1147244181, -57.8592009928, 22.0796103591, 86.3047428322, 4.30917477192, 0.861860386863, 20.5273846088, -48.1961190472};
test_label[4865] = '{20.5273846088};
test_output[4865] = '{65.7773582234};
############ END DEBUG ############*/
test_input[38928:38935] = '{32'hc0d1194a, 32'hc23375b5, 32'h3e91495f, 32'h41b78474, 32'hc251efd7, 32'hc21f6a4f, 32'hc02bc3ad, 32'h4120552e};
test_label[4866] = '{32'hc251efd7};
test_output[4866] = '{32'h4296d909};
/*############ DEBUG ############
test_input[38928:38935] = '{-6.53433686554, -44.8649475241, 0.28376290338, 22.9396740223, -52.4842179531, -39.85381573, -2.68381799949, 10.0207962583};
test_label[4866] = '{-52.4842179531};
test_output[4866] = '{75.4238944268};
############ END DEBUG ############*/
test_input[38936:38943] = '{32'h4221b0ac, 32'hc264519c, 32'hc2c0f29d, 32'h41f0bbcc, 32'hc298a9f6, 32'h428039a5, 32'hc2a0f155, 32'h428a924e};
test_label[4867] = '{32'hc2a0f155};
test_output[4867] = '{32'h4315c344};
/*############ DEBUG ############
test_input[38936:38943] = '{40.4225327959, -57.0796985148, -96.4738534577, 30.0916968772, -76.3319540548, 64.1125855372, -80.4713522646, 69.2857494914};
test_label[4867] = '{-80.4713522646};
test_output[4867] = '{149.762752373};
############ END DEBUG ############*/
test_input[38944:38951] = '{32'h423135eb, 32'hc2bea124, 32'h42a6cc3c, 32'h42b4da61, 32'h41b10a97, 32'h412db252, 32'hc2747473, 32'hc2295bcc};
test_label[4868] = '{32'h423135eb};
test_output[4868] = '{32'h42387fbf};
/*############ DEBUG ############
test_input[38944:38951] = '{44.3026549865, -95.3147261874, 83.3988962349, 90.4265187196, 22.130169927, 10.8560356398, -61.1137184695, -42.3396435659};
test_label[4868] = '{44.3026549865};
test_output[4868] = '{46.1247503781};
############ END DEBUG ############*/
test_input[38952:38959] = '{32'hc257a92f, 32'hc21fcc00, 32'hc2808996, 32'hc1c72881, 32'h4250452e, 32'hc2a84cee, 32'h426308a3, 32'hc2aa523f};
test_label[4869] = '{32'hc2aa523f};
test_output[4869] = '{32'h430ded9f};
/*############ DEBUG ############
test_input[38952:38959] = '{-53.9152202193, -39.9492197583, -64.2687231851, -24.8947768075, 52.0675592133, -84.1502534412, 56.7584341565, -85.1606364443};
test_label[4869] = '{-85.1606364443};
test_output[4869] = '{141.928207385};
############ END DEBUG ############*/
test_input[38960:38967] = '{32'h42acec29, 32'hc26cfcde, 32'hc2af8c88, 32'hc12e8212, 32'h4237a35c, 32'hc190fdbb, 32'h427fab49, 32'hc27a2621};
test_label[4870] = '{32'h427fab49};
test_output[4870] = '{32'h41b45a13};
/*############ DEBUG ############
test_input[38960:38967] = '{86.4612519883, -59.2469414956, -87.7744724018, -10.9067552765, 45.909530089, -18.1238913941, 63.9172709158, -62.5372350166};
test_label[4870] = '{63.9172709158};
test_output[4870] = '{22.5439810727};
############ END DEBUG ############*/
test_input[38968:38975] = '{32'hc1da2b10, 32'h41eb8d78, 32'h41a50f3e, 32'h404062e3, 32'hc25a7378, 32'h42c723d5, 32'hc2858ec0, 32'h426eb887};
test_label[4871] = '{32'h42c723d5};
test_output[4871] = '{32'h80000000};
/*############ DEBUG ############
test_input[38968:38975] = '{-27.2710275508, 29.4440759731, 20.6324431082, 3.00603557992, -54.6127633879, 99.5699824363, -66.7788117676, 59.680201432};
test_label[4871] = '{99.5699824363};
test_output[4871] = '{-0.0};
############ END DEBUG ############*/
test_input[38976:38983] = '{32'hc0265132, 32'hc28416e5, 32'hc221dcaf, 32'hc2bd23e1, 32'hc238c17a, 32'hc17b9bc6, 32'hc26132bd, 32'hbe6b3cb5};
test_label[4872] = '{32'hc0265132};
test_output[4872] = '{32'h401d5700};
/*############ DEBUG ############
test_input[38976:38983] = '{-2.59870570119, -66.0447176179, -40.4655128771, -94.5700735854, -46.1889406992, -15.7255307792, -56.2995481749, -0.229723773045};
test_label[4872] = '{-2.59870570119};
test_output[4872] = '{2.4584351084};
############ END DEBUG ############*/
test_input[38984:38991] = '{32'h429ee363, 32'hc2b6c543, 32'h42a38d03, 32'h4255565d, 32'h421c26ae, 32'h4121593b, 32'h42b556ec, 32'h42088c55};
test_label[4873] = '{32'h429ee363};
test_output[4873] = '{32'h41339ce7};
/*############ DEBUG ############
test_input[38984:38991] = '{79.4441157257, -91.3852742965, 81.7754106142, 53.3343380459, 39.0377729138, 10.084284432, 90.6697713492, 34.1370431414};
test_label[4873] = '{79.4441157257};
test_output[4873] = '{11.2258061002};
############ END DEBUG ############*/
test_input[38992:38999] = '{32'h41824ff8, 32'h42a0cc95, 32'h428bb410, 32'h4180dd34, 32'h41df7ac2, 32'hc2428fe3, 32'hc2bf4bee, 32'hc2c011d2};
test_label[4874] = '{32'h4180dd34};
test_output[4874] = '{32'h4280954c};
/*############ DEBUG ############
test_input[38992:38999] = '{16.289046942, 80.3995765677, 69.8516808157, 16.1080087962, 27.9349409367, -48.6405131426, -95.6482974023, -96.0348078228};
test_label[4874] = '{16.1080087962};
test_output[4874] = '{64.2915940199};
############ END DEBUG ############*/
test_input[39000:39007] = '{32'hc1f58250, 32'h42c43781, 32'h425af049, 32'hc17054b7, 32'h428de5cb, 32'hc12ccddc, 32'h40d792d4, 32'h42bb8572};
test_label[4875] = '{32'h425af049};
test_output[4875] = '{32'h422d8be3};
/*############ DEBUG ############
test_input[39000:39007] = '{-30.6886283471, 98.1084056734, 54.7346518837, -15.0206820241, 70.9488146939, -10.8002586216, 6.73667320631, 93.7606371169};
test_label[4875] = '{54.7346518837};
test_output[4875] = '{43.3866064843};
############ END DEBUG ############*/
test_input[39008:39015] = '{32'h42597d3e, 32'h4199ab13, 32'hc0ec61d4, 32'h42ab4184, 32'h41a891db, 32'h406f733c, 32'h429f7f60, 32'hc283e53d};
test_label[4876] = '{32'h429f7f60};
test_output[4876] = '{32'h40bc3923};
/*############ DEBUG ############
test_input[39008:39015] = '{54.3723062176, 19.2085329236, -7.38694173225, 85.6279601699, 21.0712179793, 3.74140842572, 79.7487787539, -65.9477289135};
test_label[4876] = '{79.7487787539};
test_output[4876] = '{5.88197458547};
############ END DEBUG ############*/
test_input[39016:39023] = '{32'h42719057, 32'h42555c34, 32'hc214af8c, 32'h40c425ab, 32'hc1995fdb, 32'h42c50bf4, 32'hc1c857dd, 32'h4218e79a};
test_label[4877] = '{32'h42719057};
test_output[4877] = '{32'h42188791};
/*############ DEBUG ############
test_input[39016:39023] = '{60.3909555, 53.3400414715, -37.1714309782, 6.12959834369, -19.1718053079, 98.5233447812, -25.0429028591, 38.2261740276};
test_label[4877] = '{60.3909555};
test_output[4877] = '{38.1323892812};
############ END DEBUG ############*/
test_input[39024:39031] = '{32'hc2a1e444, 32'hc20915d7, 32'h409c03f9, 32'h42141bd4, 32'hc2989fa2, 32'h4192aa16, 32'hbf467f37, 32'hc1768d3d};
test_label[4878] = '{32'hc1768d3d};
test_output[4878] = '{32'h4251bf23};
/*############ DEBUG ############
test_input[39024:39031] = '{-80.9458310847, -34.2713265221, 4.87548512741, 37.027175565, -76.3117841331, 18.3330495677, -0.77537862016, -15.4094818226};
test_label[4878] = '{-15.4094818226};
test_output[4878] = '{52.4366573952};
############ END DEBUG ############*/
test_input[39032:39039] = '{32'hc2c4ee9b, 32'h3ff97a98, 32'h42a4ed0a, 32'hc29ac5d1, 32'h42bd3ddf, 32'hc2b9e924, 32'hc2b4576c, 32'h422f8a43};
test_label[4879] = '{32'hc2b9e924};
test_output[4879] = '{32'h433b9382};
/*############ DEBUG ############
test_input[39032:39039] = '{-98.4660244668, 1.94905374446, 82.4629634246, -77.3863622549, 94.6208413601, -92.9553526141, -90.1707495247, 43.8850194567};
test_label[4879] = '{-92.9553526141};
test_output[4879] = '{187.576199221};
############ END DEBUG ############*/
test_input[39040:39047] = '{32'h428bac5f, 32'hc1c6fc57, 32'hc266e3f7, 32'h423a2f26, 32'h42a4224d, 32'hc21a0eff, 32'h41e2fd29, 32'h4237b794};
test_label[4880] = '{32'h423a2f26};
test_output[4880] = '{32'h420e1576};
/*############ DEBUG ############
test_input[39040:39047] = '{69.8366592071, -24.873213608, -57.7226223232, 46.5460420739, 82.0669940225, -38.5146446158, 28.373612405, 45.929276684};
test_label[4880] = '{46.5460420739};
test_output[4880] = '{35.5209568287};
############ END DEBUG ############*/
test_input[39048:39055] = '{32'hbfe68e80, 32'h400e3497, 32'h41c368ba, 32'h4285d330, 32'h423b1bc9, 32'h42ada884, 32'h419c7d7c, 32'hc2106d33};
test_label[4881] = '{32'hc2106d33};
test_output[4881] = '{32'h42f5df1e};
/*############ DEBUG ############
test_input[39048:39055] = '{-1.80122379326, 2.2219597408, 24.4261364891, 66.9124719738, 46.7771333578, 86.8291344735, 19.561272477, -36.1066408601};
test_label[4881] = '{-36.1066408601};
test_output[4881] = '{122.935775336};
############ END DEBUG ############*/
test_input[39056:39063] = '{32'h42393000, 32'hc1f4a070, 32'hc1b0256a, 32'hc1507b91, 32'hc2a47dc5, 32'hc0246545, 32'h4096fc89, 32'h42c65f20};
test_label[4882] = '{32'h4096fc89};
test_output[4882] = '{32'h42bcef58};
/*############ DEBUG ############
test_input[39056:39063] = '{46.2968764549, -30.5783377699, -22.018268606, -13.030167385, -82.2456452205, -2.56868107506, 4.71832726459, 99.1857948173};
test_label[4882] = '{4.71832726459};
test_output[4882] = '{94.4674675527};
############ END DEBUG ############*/
test_input[39064:39071] = '{32'h41ec95b9, 32'h424c2a5b, 32'h41b7bd00, 32'hc21a1177, 32'hc2b8a4f3, 32'hc1a33cc0, 32'hc0ed0139, 32'hc15c7d27};
test_label[4883] = '{32'hc0ed0139};
test_output[4883] = '{32'h4269ca82};
/*############ DEBUG ############
test_input[39064:39071] = '{29.5731070345, 51.0413619546, 22.967284605, -38.5170537643, -92.322163576, -20.4046622598, -7.40639904324, -13.7805549673};
test_label[4883] = '{-7.40639904324};
test_output[4883] = '{58.4477609983};
############ END DEBUG ############*/
test_input[39072:39079] = '{32'h4193c280, 32'hc19e4750, 32'hc09a743f, 32'h419c26e5, 32'hc26a56b6, 32'hc2bc498d, 32'hc2ad1b20, 32'h4285d073};
test_label[4884] = '{32'hc26a56b6};
test_output[4884] = '{32'h42fafbce};
/*############ DEBUG ############
test_input[39072:39079] = '{18.4699701186, -19.7848205325, -4.82669000883, 19.5189921659, -58.5846787916, -94.1436533304, -86.5529766209, 66.9071281964};
test_label[4884] = '{-58.5846787916};
test_output[4884] = '{125.491806988};
############ END DEBUG ############*/
test_input[39080:39087] = '{32'h41900db2, 32'h4186e2a6, 32'h421ec29d, 32'h41a602d9, 32'h42a18de9, 32'h416bb085, 32'hc2b7e52c, 32'h41776ecb};
test_label[4885] = '{32'h416bb085};
test_output[4885] = '{32'h428417d9};
/*############ DEBUG ############
test_input[39080:39087] = '{18.0066880724, 16.8606682176, 39.6900536883, 20.7513906053, 80.7771713567, 14.7305954711, -91.9475993248, 15.4645486525};
test_label[4885] = '{14.7305954711};
test_output[4885] = '{66.0465758856};
############ END DEBUG ############*/
test_input[39088:39095] = '{32'hc2029d35, 32'h420b921e, 32'h411358b7, 32'h41997006, 32'h42b9ace6, 32'hc27a73c3, 32'h420f7f16, 32'hc2c69ca0};
test_label[4886] = '{32'h420b921e};
test_output[4886] = '{32'h4267c7ad};
/*############ DEBUG ############
test_input[39088:39095] = '{-32.6535229007, 34.8926925188, 9.20915914306, 19.1796989733, 92.8376885974, -62.6130470529, 35.8741091491, -99.3059101816};
test_label[4886] = '{34.8926925188};
test_output[4886] = '{57.9449960786};
############ END DEBUG ############*/
test_input[39096:39103] = '{32'h42c72a41, 32'hc1c0e52b, 32'hc27f9b2f, 32'hc120af72, 32'h42892177, 32'h42c137f7, 32'h42b409af, 32'h412f8e1e};
test_label[4887] = '{32'h412f8e1e};
test_output[4887] = '{32'h42b1520f};
/*############ DEBUG ############
test_input[39096:39103] = '{99.582524947, -24.1118984851, -63.9015469474, -10.0428332414, 68.5653629416, 96.6093076744, 90.0189145162, 10.9721963843};
test_label[4887] = '{10.9721963843};
test_output[4887] = '{88.6602692624};
############ END DEBUG ############*/
test_input[39104:39111] = '{32'hc2c19904, 32'h428a5608, 32'hc080fde5, 32'h42a901df, 32'h42b34f28, 32'hc26ea4ce, 32'h42bb53ec, 32'h41694ac4};
test_label[4888] = '{32'h42b34f28};
test_output[4888] = '{32'h4080e06f};
/*############ DEBUG ############
test_input[39104:39111] = '{-96.7988564523, 69.1680293548, -4.03099307885, 84.5036552648, 89.6545989379, -59.6609415101, 93.6639089073, 14.5807531148};
test_label[4888] = '{89.6545989379};
test_output[4888] = '{4.02739646657};
############ END DEBUG ############*/
test_input[39112:39119] = '{32'hc22b62e5, 32'h41c88ab5, 32'hc293814e, 32'hc205355e, 32'h3fe79fa3, 32'hc17288d4, 32'h3f8e23c9, 32'hc11bda27};
test_label[4889] = '{32'hc17288d4};
test_output[4889] = '{32'h4220e78f};
/*############ DEBUG ############
test_input[39112:39119] = '{-42.8465761774, 25.0677276878, -73.7525463704, -33.3021162586, 1.80955923405, -15.1584049741, 1.11046704039, -9.74075967207};
test_label[4889] = '{-15.1584049741};
test_output[4889] = '{40.226132662};
############ END DEBUG ############*/
test_input[39120:39127] = '{32'h42c31139, 32'hc199e9eb, 32'h4254b754, 32'hc224e895, 32'h40942d3d, 32'hc1a67410, 32'hc2b4d4ce, 32'h423d5125};
test_label[4890] = '{32'hc224e895};
test_output[4890] = '{32'h430ac2c2};
/*############ DEBUG ############
test_input[39120:39127] = '{97.533638766, -19.2392183827, 53.1790328395, -41.2271297873, 4.63052212659, -20.8066705137, -90.4156349465, 47.329244146};
test_label[4890] = '{-41.2271297873};
test_output[4890] = '{138.760768553};
############ END DEBUG ############*/
test_input[39128:39135] = '{32'hc27e14cf, 32'h42a31752, 32'hc26af36e, 32'hc2a6e303, 32'hc2b55d10, 32'h424ebbc0, 32'h4126e892, 32'hc2c0f4d2};
test_label[4891] = '{32'hc27e14cf};
test_output[4891] = '{32'h431110dd};
/*############ DEBUG ############
test_input[39128:39135] = '{-63.520322546, 81.5455469045, -58.737723125, -83.4433792742, -90.6817640237, 51.6833511773, 10.4317795169, -96.4781658972};
test_label[4891] = '{-63.520322546};
test_output[4891] = '{145.065869451};
############ END DEBUG ############*/
test_input[39136:39143] = '{32'h40b4ee51, 32'h42b32fa4, 32'h42136847, 32'hc2953e10, 32'h421c3a95, 32'h42883137, 32'h4253a114, 32'hc20c0c7a};
test_label[4892] = '{32'h42b32fa4};
test_output[4892] = '{32'h2ffd9d24};
/*############ DEBUG ############
test_input[39136:39143] = '{5.65409132463, 89.5930481471, 36.8518315933, -74.6212189311, 39.0572100146, 68.096120763, 52.9073028741, -35.0121833947};
test_label[4892] = '{89.5930481471};
test_output[4892] = '{4.61320870499e-10};
############ END DEBUG ############*/
test_input[39144:39151] = '{32'h40e30f61, 32'hc0fe438f, 32'h4104161d, 32'hc2a5caed, 32'h3dc3b274, 32'hc0550a05, 32'h40ae6f34, 32'h42b17c22};
test_label[4893] = '{32'h40e30f61};
test_output[4893] = '{32'h42a34b2c};
/*############ DEBUG ############
test_input[39144:39151] = '{7.09562741948, -7.94574697896, 8.2553985301, -82.8963367396, 0.0955552135984, -3.32873653836, 5.45107477575, 88.7424450846};
test_label[4893] = '{7.09562741948};
test_output[4893] = '{81.6468176651};
############ END DEBUG ############*/
test_input[39152:39159] = '{32'h428f6e0a, 32'h41655179, 32'h427eb255, 32'hc2775047, 32'hc2825708, 32'h423c9ae4, 32'hc27acecc, 32'hc23344d1};
test_label[4894] = '{32'hc2775047};
test_output[4894] = '{32'h43058b2c};
/*############ DEBUG ############
test_input[39152:39159] = '{71.7149213801, 14.332390498, 63.6741541001, -61.8283954189, -65.169983565, 47.1512619411, -62.7019500899, -44.817203813};
test_label[4894] = '{-61.8283954189};
test_output[4894] = '{133.543638809};
############ END DEBUG ############*/
test_input[39160:39167] = '{32'hc1501267, 32'h41ef71d0, 32'h40aeb6a0, 32'h42380d4f, 32'h42ade397, 32'h425f16ea, 32'h42704fcd, 32'h424a6429};
test_label[4895] = '{32'h425f16ea};
test_output[4895] = '{32'h41f9608a};
/*############ DEBUG ############
test_input[39160:39167] = '{-13.0044923239, 29.9305730552, 5.459792899, 46.0129949724, 86.9445129499, 55.7723756363, 60.077930764, 50.5978126962};
test_label[4895] = '{55.7723756363};
test_output[4895] = '{31.1721373136};
############ END DEBUG ############*/
test_input[39168:39175] = '{32'h411ee6d5, 32'hc1c445fa, 32'h40a30fe8, 32'h417674fb, 32'h4247fa4c, 32'hc2a36573, 32'h40ea9be0, 32'hc0fc94be};
test_label[4896] = '{32'h411ee6d5};
test_output[4896] = '{32'h42204097};
/*############ DEBUG ############
test_input[39168:39175] = '{9.93135573657, -24.5341679969, 5.09569174519, 15.4035600604, 49.9944299295, -81.6981428116, 7.3315277376, -7.89315697075};
test_label[4896] = '{9.93135573657};
test_output[4896] = '{40.0630741929};
############ END DEBUG ############*/
test_input[39176:39183] = '{32'h429788ff, 32'hc2b2deb5, 32'h4101bf56, 32'hc143cb47, 32'hbfff248a, 32'h429aa59c, 32'h41855ff9, 32'h41cfd06d};
test_label[4897] = '{32'hc2b2deb5};
test_output[4897] = '{32'h4326f32b};
/*############ DEBUG ############
test_input[39176:39183] = '{75.767571428, -89.4349717465, 8.10921313468, -12.2371279549, -1.993302557, 77.3234552945, 16.6718624635, 25.9767707629};
test_label[4897] = '{-89.4349717465};
test_output[4897] = '{166.949875819};
############ END DEBUG ############*/
test_input[39184:39191] = '{32'h4299dd77, 32'hc1a5cffa, 32'hc2929a48, 32'h429de266, 32'h426c6306, 32'hc180952f, 32'hc1cd97af, 32'hc2a48d24};
test_label[4898] = '{32'hc180952f};
test_output[4898] = '{32'h42be4819};
/*############ DEBUG ############
test_input[39184:39191] = '{76.9325476621, -20.726551409, -73.3013276017, 78.9421866425, 59.0967030808, -16.0728426708, -25.6990638162, -82.2756640904};
test_label[4898] = '{-16.0728426708};
test_output[4898] = '{95.1408131974};
############ END DEBUG ############*/
test_input[39192:39199] = '{32'hc208f5ed, 32'h42a46d8c, 32'h422975cb, 32'hc28ecf74, 32'h42a7dcae, 32'h424bc163, 32'h423eb295, 32'h4051b9ca};
test_label[4899] = '{32'h423eb295};
test_output[4899] = '{32'h4211afea};
/*############ DEBUG ############
test_input[39192:39199] = '{-34.2401613711, 82.2139567118, 42.365032179, -71.4051812029, 83.9310176025, 50.9388539218, 47.6743960318, 3.27696471521};
test_label[4899] = '{47.6743960318};
test_output[4899] = '{36.4217912184};
############ END DEBUG ############*/
test_input[39200:39207] = '{32'hc26f9bcc, 32'hc19f7fdb, 32'h42ab37df, 32'hc230e062, 32'h41f83f7b, 32'hc13b36d9, 32'hc01f1300, 32'hc28cf692};
test_label[4900] = '{32'hc19f7fdb};
test_output[4900] = '{32'h42d317d6};
/*############ DEBUG ############
test_input[39200:39207] = '{-59.9021442002, -19.9374302928, 85.6091257109, -44.2191232115, 31.0309958772, -11.7008906759, -2.4855346257, -70.4815862814};
test_label[4900] = '{-19.9374302928};
test_output[4900] = '{105.546556004};
############ END DEBUG ############*/
test_input[39208:39215] = '{32'hc2b165d8, 32'h42aafe5f, 32'hc1e737b9, 32'h41c67d79, 32'hc2a67f3a, 32'h4295a5c1, 32'hc2a28788, 32'h41c2c7ce};
test_label[4901] = '{32'h42aafe5f};
test_output[4901] = '{32'h37c24779};
/*############ DEBUG ############
test_input[39208:39215] = '{-88.6989099366, 85.4968147933, -28.9022076549, 24.8112664104, -83.2484868915, 74.8237374815, -81.2647056711, 24.347559991};
test_label[4901] = '{85.4968147933};
test_output[4901] = '{2.31598845108e-05};
############ END DEBUG ############*/
test_input[39216:39223] = '{32'h40bb0ba4, 32'h41ad949e, 32'hc28e49f1, 32'h4158fa8f, 32'h428012ff, 32'hc2930e7f, 32'h42963bbe, 32'h41a0007b};
test_label[4902] = '{32'h41ad949e};
test_output[4902] = '{32'h4255ad30};
/*############ DEBUG ############
test_input[39216:39223] = '{5.84517075361, 21.6975674014, -71.1444153793, 13.5611718706, 64.0371030029, -73.5283123482, 75.1166810936, 20.0002336979};
test_label[4902] = '{21.6975674014};
test_output[4902] = '{53.4191291163};
############ END DEBUG ############*/
test_input[39224:39231] = '{32'h41aca6c2, 32'h421b5d14, 32'h3f668424, 32'hbfa12aa4, 32'h4217d270, 32'hc13f2672, 32'h41e4b5c1, 32'h42b1fa29};
test_label[4903] = '{32'h41e4b5c1};
test_output[4903] = '{32'h42719972};
/*############ DEBUG ############
test_input[39224:39231] = '{21.5814249444, 38.8408962156, 0.900453830406, -1.259113768, 37.9555071672, -11.946885784, 28.5887468001, 88.9885963745};
test_label[4903] = '{28.5887468001};
test_output[4903] = '{60.3998495744};
############ END DEBUG ############*/
test_input[39232:39239] = '{32'h4266c8ae, 32'h429f622c, 32'hc2a6eca5, 32'h40feed75, 32'hc2677a91, 32'hc10cbbff, 32'h40d5a2ba, 32'h428cb983};
test_label[4904] = '{32'h428cb983};
test_output[4904] = '{32'h411545a4};
/*############ DEBUG ############
test_input[39232:39239] = '{57.6959766931, 79.6917433093, -83.4621959621, 7.96648642735, -57.8696933235, -8.79589702451, 6.67611410338, 70.3623299165};
test_label[4904] = '{70.3623299165};
test_output[4904] = '{9.32950216347};
############ END DEBUG ############*/
test_input[39240:39247] = '{32'hc15afd0a, 32'h42aa57ed, 32'hc12ae49a, 32'hc1e1703b, 32'hc280bcdc, 32'h40ccdfa3, 32'hc2afde26, 32'h41faacfc};
test_label[4905] = '{32'hc2afde26};
test_output[4905] = '{32'h432d1b0a};
/*############ DEBUG ############
test_input[39240:39247] = '{-13.6867770546, 85.1717336876, -10.6808112253, -28.17979958, -64.3688664407, 6.40229939892, -87.9338818914, 31.3344650409};
test_label[4905] = '{-87.9338818914};
test_output[4905] = '{173.105615579};
############ END DEBUG ############*/
test_input[39248:39255] = '{32'hc29d4b20, 32'hc29ea318, 32'hc1aeacb5, 32'h42b4a610, 32'hc2c55568, 32'h419dd1d9, 32'h42b353f2, 32'h42abf57b};
test_label[4906] = '{32'hc2c55568};
test_output[4906] = '{32'h433d6a8a};
/*############ DEBUG ############
test_input[39248:39255] = '{-78.646730921, -79.3185401037, -21.8343295158, 90.3243437952, -98.6668081111, 19.7274656146, 89.6639518976, 85.9794517045};
test_label[4906] = '{-98.6668081111};
test_output[4906] = '{189.416172375};
############ END DEBUG ############*/
test_input[39256:39263] = '{32'hc10fa7dc, 32'hc2aed654, 32'h41f95484, 32'hc1ff08b8, 32'hc2819a84, 32'hc0cfaf41, 32'hc29147fc, 32'hc23b95f0};
test_label[4907] = '{32'hc10fa7dc};
test_output[4907] = '{32'h42209439};
/*############ DEBUG ############
test_input[39256:39263] = '{-8.97848097498, -87.4186105785, 31.1662679466, -31.879258155, -64.8017853761, -6.49014319596, -72.6405921412, -46.8964225607};
test_label[4907] = '{-8.97848097498};
test_output[4907] = '{40.1447489216};
############ END DEBUG ############*/
test_input[39264:39271] = '{32'hc2ac6ea0, 32'h41900416, 32'h42b5519b, 32'h41aa9bd0, 32'h42c1fafd, 32'h421e5246, 32'hc0f3a97b, 32'hc207da07};
test_label[4908] = '{32'hc207da07};
test_output[4908] = '{32'h4302f475};
/*############ DEBUG ############
test_input[39264:39271] = '{-86.2160654597, 18.0019950464, 90.6593871516, 21.3260795945, 96.9902114263, 39.5803464735, -7.61443861406, -33.9629172356};
test_label[4908] = '{-33.9629172356};
test_output[4908] = '{130.954907644};
############ END DEBUG ############*/
test_input[39272:39279] = '{32'hc29d6c24, 32'hc2bd51fc, 32'h4281687c, 32'hc29984ad, 32'h4257ac00, 32'h42a0a1c1, 32'hc1e7e170, 32'h40db27e1};
test_label[4909] = '{32'hc29d6c24};
test_output[4909] = '{32'h431f06f3};
/*############ DEBUG ############
test_input[39272:39279] = '{-78.7112100027, -94.6601280674, 64.7040701393, -76.7591302678, 53.9179700247, 80.3159290782, -28.9850762845, 6.84861780097};
test_label[4909] = '{-78.7112100027};
test_output[4909] = '{159.027139247};
############ END DEBUG ############*/
test_input[39280:39287] = '{32'h42598c2b, 32'h429fa44d, 32'h424a6797, 32'h411c18c6, 32'hc2a01bcb, 32'hc26f411a, 32'hc177a45a, 32'hc2a88e4b};
test_label[4910] = '{32'hc2a88e4b};
test_output[4910] = '{32'h4324194c};
/*############ DEBUG ############
test_input[39280:39287] = '{54.386882604, 79.8209002882, 50.6011606551, 9.75604826524, -80.0542803522, -59.8135763303, -15.4776251686, -84.2779187126};
test_label[4910] = '{-84.2779187126};
test_output[4910] = '{164.098819001};
############ END DEBUG ############*/
test_input[39288:39295] = '{32'h413fe82a, 32'hc2b6adb9, 32'h42b82854, 32'h42548728, 32'h41ffd89c, 32'h421f0fd9, 32'h41759f66, 32'hc2c13a2f};
test_label[4911] = '{32'hc2b6adb9};
test_output[4911] = '{32'h43376b07};
/*############ DEBUG ############
test_input[39288:39295] = '{11.9941806086, -91.339298769, 92.0787695691, 53.1319888473, 31.9807666452, 39.7654747462, 15.3514157225, -96.6136368957};
test_label[4911] = '{-91.339298769};
test_output[4911] = '{183.418068338};
############ END DEBUG ############*/
test_input[39296:39303] = '{32'hc1b6800d, 32'hc20c944b, 32'hc28d31fc, 32'h41f17380, 32'h42790416, 32'h403f1945, 32'h411961bb, 32'h42b1da8e};
test_label[4912] = '{32'h411961bb};
test_output[4912] = '{32'h429eae56};
/*############ DEBUG ############
test_input[39296:39303] = '{-22.8125242681, -35.1448165618, -70.5976242539, 30.1813959797, 62.2539890352, 2.98591729846, 9.58636022867, 88.9268631713};
test_label[4912] = '{9.58636022867};
test_output[4912] = '{79.3405029427};
############ END DEBUG ############*/
test_input[39304:39311] = '{32'hc28fa847, 32'hc1c43fb4, 32'h42038de4, 32'h42af4806, 32'hc2853cf0, 32'hc226071f, 32'hc252344b, 32'hc28ed00a};
test_label[4913] = '{32'hc2853cf0};
test_output[4913] = '{32'h431a427b};
/*############ DEBUG ############
test_input[39304:39311] = '{-71.8286674261, -24.5311054676, 32.8885649288, 87.6406705857, -66.6190178876, -41.5069552079, -52.5510685317, -71.4063261641};
test_label[4913] = '{-66.6190178876};
test_output[4913] = '{154.259688473};
############ END DEBUG ############*/
test_input[39312:39319] = '{32'hc287e8fe, 32'h42697671, 32'hc21d0cf9, 32'h413c1907, 32'hc2b7f0e7, 32'h429b3455, 32'hc2b5c939, 32'hc21c01a7};
test_label[4914] = '{32'hc21d0cf9};
test_output[4914] = '{32'h42e9bad2};
/*############ DEBUG ############
test_input[39312:39319] = '{-67.9550614312, 58.365663889, -39.2626669441, 11.7561105497, -91.9705116926, 77.6022130704, -90.8930138051, -39.0016139185};
test_label[4914] = '{-39.2626669441};
test_output[4914] = '{116.864880019};
############ END DEBUG ############*/
test_input[39320:39327] = '{32'h42905060, 32'hc19aa77a, 32'hc1c2ad92, 32'h414568dc, 32'hc0b5eaa8, 32'h41405b16, 32'hc26fb698, 32'h42b41ee4};
test_label[4915] = '{32'h42905060};
test_output[4915] = '{32'h418f3a0c};
/*############ DEBUG ############
test_input[39320:39327] = '{72.1569858546, -19.3317751969, -24.3347519498, 12.3381007823, -5.6848947091, 12.0222374948, -59.9283153883, 90.0603299566};
test_label[4915] = '{72.1569858546};
test_output[4915] = '{17.9033441187};
############ END DEBUG ############*/
test_input[39328:39335] = '{32'h42196487, 32'hc28a8b12, 32'hc109e282, 32'hc0627f4d, 32'h42a06278, 32'h42bed937, 32'hc259a809, 32'hc2b27e31};
test_label[4916] = '{32'h42a06278};
test_output[4916] = '{32'h4173b5fc};
/*############ DEBUG ############
test_input[39328:39335] = '{38.3481715731, -69.2716253377, -8.61779964289, -3.53901990314, 80.1923209659, 95.4242506916, -54.4140961699, -89.2464670377};
test_label[4916] = '{80.1923209659};
test_output[4916] = '{15.2319299683};
############ END DEBUG ############*/
test_input[39336:39343] = '{32'hc277c4ed, 32'hc0bd2557, 32'hc29c98cb, 32'hc1e329f3, 32'h417ce956, 32'h42a7b66d, 32'hc1a2c128, 32'hc0a0e06e};
test_label[4917] = '{32'h417ce956};
test_output[4917] = '{32'h42881942};
/*############ DEBUG ############
test_input[39336:39343] = '{-61.9423084418, -5.9108081454, -78.2984273287, -28.3954822548, 15.8069672413, 83.8563000803, -20.3443138665, -5.02739605947};
test_label[4917] = '{15.8069672413};
test_output[4917] = '{68.049332839};
############ END DEBUG ############*/
test_input[39344:39351] = '{32'hc28ad32b, 32'hc1a185bb, 32'h42b50f4e, 32'hc255228b, 32'h4271003f, 32'h42b3db28, 32'hc20de92b, 32'h41850d29};
test_label[4918] = '{32'h42b3db28};
test_output[4918] = '{32'h3f84f37e};
/*############ DEBUG ############
test_input[39344:39351] = '{-69.4124359481, -20.1902976087, 90.5298899234, -53.2837327081, 60.2502407316, 89.9280430925, -35.4777030988, 16.6314256055};
test_label[4918] = '{89.9280430925};
test_output[4918] = '{1.03868075858};
############ END DEBUG ############*/
test_input[39352:39359] = '{32'h41f2c0b9, 32'h428a7cfd, 32'h41edba52, 32'hc1ad522d, 32'hc2b7876b, 32'h41d96cd3, 32'hc08c12f5, 32'h42915e9f};
test_label[4919] = '{32'h41edba52};
test_output[4919] = '{32'h422c0061};
/*############ DEBUG ############
test_input[39352:39359] = '{30.3441026225, 69.2441152522, 29.7159760667, -21.6651244362, -91.7644892241, 27.1781371673, -4.3773140257, 72.6848075631};
test_label[4919] = '{29.7159760667};
test_output[4919] = '{43.0003713393};
############ END DEBUG ############*/
test_input[39360:39367] = '{32'h429ce936, 32'hc2ba48fb, 32'hc227f688, 32'h408320c9, 32'h4225c154, 32'hc2291736, 32'h42371163, 32'h426d8199};
test_label[4920] = '{32'h4225c154};
test_output[4920] = '{32'h42141118};
/*############ DEBUG ############
test_input[39360:39367] = '{78.4554888023, -93.1425413784, -41.990751293, 4.09775226366, 41.4387952919, -42.2726664828, 45.7669805534, 59.3765597406};
test_label[4920] = '{41.4387952919};
test_output[4920] = '{37.0166935156};
############ END DEBUG ############*/
test_input[39368:39375] = '{32'hc28a5934, 32'h42bfba01, 32'hc2c2a082, 32'h42431297, 32'hc2bea548, 32'hc14eda6f, 32'hc2b791ed, 32'hc2333c79};
test_label[4921] = '{32'hc28a5934};
test_output[4921] = '{32'h4325099b};
/*############ DEBUG ############
test_input[39368:39375] = '{-69.1742279912, 95.8632899208, -97.313494847, 48.7681554206, -95.3228132542, -12.9283282744, -91.7850093663, -44.8090539637};
test_label[4921] = '{-69.1742279912};
test_output[4921] = '{165.037517912};
############ END DEBUG ############*/
test_input[39376:39383] = '{32'h42bd82aa, 32'h428e6017, 32'hc2aca12e, 32'hc2adaefb, 32'h429549c5, 32'hc264d1b8, 32'h426ca3f5, 32'hc28ff747};
test_label[4922] = '{32'hc264d1b8};
test_output[4922] = '{32'h4317f5c3};
/*############ DEBUG ############
test_input[39376:39383] = '{94.7552020374, 71.1876752532, -86.3148071478, -86.8417562437, 74.6440848982, -57.2048035306, 59.1601151862, -71.9829646154};
test_label[4922] = '{-57.2048035306};
test_output[4922] = '{151.96000557};
############ END DEBUG ############*/
test_input[39384:39391] = '{32'hc22ef2e9, 32'hbf026d38, 32'hc295fd76, 32'hc29734e2, 32'hc1b613d6, 32'h412f0445, 32'h42983f36, 32'hc24f49db};
test_label[4923] = '{32'h412f0445};
test_output[4923] = '{32'h42825eae};
/*############ DEBUG ############
test_input[39384:39391] = '{-43.7372175599, -0.50947903683, -74.9950441141, -75.6032873195, -22.7596863127, 10.9385426277, 76.1234615039, -51.8221237116};
test_label[4923] = '{10.9385426277};
test_output[4923] = '{65.1849188762};
############ END DEBUG ############*/
test_input[39392:39399] = '{32'hc23cc535, 32'h40dbcd10, 32'h42ac914c, 32'hc2bbdcb0, 32'h40fcd47e, 32'h42bb0988, 32'hc2991df2, 32'h42ba0ae5};
test_label[4924] = '{32'hc23cc535};
test_output[4924] = '{32'h430d2fce};
/*############ DEBUG ############
test_input[39392:39399] = '{-47.1925862061, 6.86878210802, 86.2837843027, -93.9310285593, 7.90093885723, 93.5186145102, -76.5584893198, 93.0212792693};
test_label[4924] = '{-47.1925862061};
test_output[4924] = '{141.186732849};
############ END DEBUG ############*/
test_input[39400:39407] = '{32'h4098aeb0, 32'h429c7e18, 32'hc2baa523, 32'hc2116080, 32'h42a53cf9, 32'h4188f8d4, 32'h4226253c, 32'h42a66368};
test_label[4925] = '{32'h42a66368};
test_output[4925] = '{32'h3ee6e001};
/*############ DEBUG ############
test_input[39400:39407] = '{4.7713242541, 78.2462795333, -93.3225355022, -36.3442391077, 82.6190909391, 17.1214988603, 41.5363609624, 83.1941539528};
test_label[4925] = '{83.1941539528};
test_output[4925] = '{0.450927769625};
############ END DEBUG ############*/
test_input[39408:39415] = '{32'hc0893849, 32'hc247e5eb, 32'hc25068c6, 32'h425d0c36, 32'h42b42cf0, 32'hc1c72bb0, 32'hc00ade03, 32'hc16cbb1f};
test_label[4926] = '{32'hc0893849};
test_output[4926] = '{32'h42bcc074};
/*############ DEBUG ############
test_input[39408:39415] = '{-4.28812075811, -49.9745293488, -52.1023185156, 55.2619265935, 90.0877665228, -24.8963325708, -2.16980045228, -14.7956834032};
test_label[4926] = '{-4.28812075811};
test_output[4926] = '{94.3758872809};
############ END DEBUG ############*/
test_input[39416:39423] = '{32'hc1c83e7e, 32'hc21776b3, 32'hc29cbf9f, 32'h402a919d, 32'h422223be, 32'hc1e1cb67, 32'hc25b310c, 32'h42b09b7c};
test_label[4927] = '{32'h422223be};
test_output[4927] = '{32'h423f133b};
/*############ DEBUG ############
test_input[39416:39423] = '{-25.030513976, -37.8659184698, -78.3742633037, 2.66513755875, 40.5349040028, -28.2243169362, -54.7978979301, 88.3036834155};
test_label[4927] = '{40.5349040028};
test_output[4927] = '{47.7687794127};
############ END DEBUG ############*/
test_input[39424:39431] = '{32'h4284a918, 32'hc29cb09e, 32'hc247fff0, 32'hc291dd5a, 32'h429402b9, 32'hc20b0f38, 32'h4266740b, 32'h429b2b71};
test_label[4928] = '{32'hc291dd5a};
test_output[4928] = '{32'h43168b71};
/*############ DEBUG ############
test_input[39424:39431] = '{66.3302625031, -78.3449527204, -49.9999372669, -72.9323302253, 74.0053144991, -34.7648604213, 57.6133232189, 77.5848432416};
test_label[4928] = '{-72.9323302253};
test_output[4928] = '{150.544693092};
############ END DEBUG ############*/
test_input[39432:39439] = '{32'h42b413d2, 32'h4131d240, 32'hc29b56ab, 32'h4229e0ba, 32'h42455079, 32'h421d8e78, 32'h429b720d, 32'h42c75305};
test_label[4929] = '{32'h4229e0ba};
test_output[4929] = '{32'h4264c562};
/*############ DEBUG ############
test_input[39432:39439] = '{90.0387133989, 11.1138307396, -77.6692749893, 42.4694589698, 49.3285868191, 39.389131188, 77.7227579196, 99.6621484559};
test_label[4929] = '{42.4694589698};
test_output[4929] = '{57.1927556442};
############ END DEBUG ############*/
test_input[39440:39447] = '{32'h425c0649, 32'hc187f8af, 32'hc2652e07, 32'h423c3a84, 32'h42322273, 32'h426b759e, 32'h42088a64, 32'h417ba6ca};
test_label[4930] = '{32'hc187f8af};
test_output[4930] = '{32'h4297c3ac};
/*############ DEBUG ############
test_input[39440:39447] = '{55.0061378588, -16.9964269209, -57.2949469607, 47.0571433417, 44.5336418665, 58.8648617327, 34.1351479873, 15.7282197409};
test_label[4930] = '{-16.9964269209};
test_output[4930] = '{75.8821720163};
############ END DEBUG ############*/
test_input[39448:39455] = '{32'h429583a9, 32'hc2886055, 32'h4285f2b5, 32'h3e18e123, 32'hc20b8aee, 32'h417caf2f, 32'h41bfd92d, 32'h3f8525a3};
test_label[4931] = '{32'h417caf2f};
test_output[4931] = '{32'h426bdbf4};
/*############ DEBUG ############
test_input[39448:39455] = '{74.7571505277, -68.1881454125, 66.9740356115, 0.14929633067, -34.8856720706, 15.7927693734, 23.9810425006, 1.04021113864};
test_label[4931] = '{15.7927693734};
test_output[4931] = '{58.9647977796};
############ END DEBUG ############*/
test_input[39456:39463] = '{32'h42bac53f, 32'hc2498dd2, 32'hc2ae18f3, 32'hc20d9af7, 32'hbf27ef21, 32'h42a8b82f, 32'hc2bba979, 32'h4186bd90};
test_label[4932] = '{32'hc2ae18f3};
test_output[4932] = '{32'h43346f21};
/*############ DEBUG ############
test_input[39456:39463] = '{93.3852441521, -50.3884971682, -87.0487298598, -35.4013314525, -0.655992585941, 84.3597316822, -93.8310008461, 16.8425602801};
test_label[4932] = '{-87.0487298598};
test_output[4932] = '{180.434094306};
############ END DEBUG ############*/
test_input[39464:39471] = '{32'h42893ca3, 32'hc2a34ca8, 32'h42aaa679, 32'h421ed66b, 32'h411a4841, 32'h42872730, 32'h418c37c0, 32'hc29eaae3};
test_label[4933] = '{32'hc29eaae3};
test_output[4933] = '{32'h4324a8ae};
/*############ DEBUG ############
test_input[39464:39471] = '{68.6184309961, -81.6497179316, 85.3251413613, 39.7093921023, 9.64263984204, 67.5765351467, 17.5272220162, -79.3337602457};
test_label[4933] = '{-79.3337602457};
test_output[4933] = '{164.658901682};
############ END DEBUG ############*/
test_input[39472:39479] = '{32'h42b28958, 32'h41d5712e, 32'hc1a84b6c, 32'hc235caad, 32'h428368d3, 32'h424938c0, 32'hc280f943, 32'h42a7ae5b};
test_label[4934] = '{32'hc235caad};
test_output[4934] = '{32'h4306b876};
/*############ DEBUG ############
test_input[39472:39479] = '{89.2682467235, 26.6802638949, -21.0368268209, -45.4479256596, 65.7047357173, 50.3054186368, -64.4868405929, 83.8405385443};
test_label[4934] = '{-45.4479256596};
test_output[4934] = '{134.720555914};
############ END DEBUG ############*/
test_input[39480:39487] = '{32'hc2aaae02, 32'h41a6bf56, 32'h423c25d1, 32'h42c6eaa7, 32'h41ef60ef, 32'hc23dc312, 32'h41c457a4, 32'h4268bb90};
test_label[4935] = '{32'h423c25d1};
test_output[4935] = '{32'h4251af7c};
/*############ DEBUG ############
test_input[39480:39487] = '{-85.3398609012, 20.8434254518, 47.0369300356, 99.4583025961, 29.9223314673, -47.440499189, 24.5427938525, 58.1831651983};
test_label[4935] = '{47.0369300356};
test_output[4935] = '{52.4213725605};
############ END DEBUG ############*/
test_input[39488:39495] = '{32'h42af1d06, 32'h42711a3b, 32'hc1b19e55, 32'h4212a373, 32'h42b9f49c, 32'hc1e39b4a, 32'h4296839d, 32'hc2803339};
test_label[4936] = '{32'h4296839d};
test_output[4936] = '{32'h418dcd05};
/*############ DEBUG ############
test_input[39488:39495] = '{87.5566868838, 60.2756170375, -22.2023107063, 36.6596172837, 92.9777514975, -28.4508253387, 75.257056834, -64.100046685};
test_label[4936] = '{75.257056834};
test_output[4936] = '{17.7251073693};
############ END DEBUG ############*/
test_input[39496:39503] = '{32'hc2b21279, 32'h42bdb1d7, 32'hc291a45e, 32'h4229994d, 32'h41cecf99, 32'h42465cf7, 32'hc2b0307e, 32'hc2489c5d};
test_label[4937] = '{32'h42bdb1d7};
test_output[4937] = '{32'h80000000};
/*############ DEBUG ############
test_input[39496:39503] = '{-89.0360793189, 94.8473429712, -72.8210330172, 42.3997075198, 25.8513651535, 49.5907871036, -88.0947140762, -50.1527001062};
test_label[4937] = '{94.8473429712};
test_output[4937] = '{-0.0};
############ END DEBUG ############*/
test_input[39504:39511] = '{32'hc2669357, 32'h41b8e7a2, 32'hc22c9793, 32'h41b3be78, 32'hc2bf4672, 32'h4154d288, 32'hc232964a, 32'h425f3ead};
test_label[4938] = '{32'hc22c9793};
test_output[4938] = '{32'h42c5eb20};
/*############ DEBUG ############
test_input[39504:39511] = '{-57.6438868488, 23.11310204, -43.1480231367, 22.4680017661, -95.6375859467, 13.3013996282, -44.6467665898, 55.8112078991};
test_label[4938] = '{-43.1480231367};
test_output[4938] = '{98.9592310358};
############ END DEBUG ############*/
test_input[39512:39519] = '{32'hc24d04fa, 32'hc037e26c, 32'h428cfd58, 32'hc229b242, 32'h41ce25d7, 32'h42b6ca4e, 32'hc1a8d5c6, 32'hc14abc46};
test_label[4939] = '{32'hc14abc46};
test_output[4939] = '{32'h42d021d7};
/*############ DEBUG ############
test_input[39512:39519] = '{-51.2548600769, -2.87319460245, 70.4948116497, -42.4240802191, 25.7684761156, 91.3951300442, -21.1043819731, -12.6709654939};
test_label[4939] = '{-12.6709654939};
test_output[4939] = '{104.066095539};
############ END DEBUG ############*/
test_input[39520:39527] = '{32'hc11f48d5, 32'hc0ad06be, 32'h42a99813, 32'h42345f3b, 32'h41f3a002, 32'h419e3df7, 32'hc27d8469, 32'h429e47c9};
test_label[4940] = '{32'h42a99813};
test_output[4940] = '{32'h3b648f74};
/*############ DEBUG ############
test_input[39520:39527] = '{-9.95528142, -5.40707298018, 84.7970162221, 45.0929968921, 30.4531297256, 19.7802557918, -63.3793061533, 79.1402059908};
test_label[4940] = '{84.7970162221};
test_output[4940] = '{0.0034875544629};
############ END DEBUG ############*/
test_input[39528:39535] = '{32'hc197fc85, 32'hc26f5de8, 32'hc2a80d1a, 32'hc2b7913d, 32'h42be4e8e, 32'h425d4934, 32'hc22b6f14, 32'h42bc2739};
test_label[4941] = '{32'hc197fc85};
test_output[4941] = '{32'h42e4e3ca};
/*############ DEBUG ############
test_input[39528:39535] = '{-18.9983008231, -59.8417050191, -84.0255923615, -91.783669677, 95.1534275262, 55.3214874647, -42.8584766007, 94.0766035776};
test_label[4941] = '{-18.9983008231};
test_output[4941] = '{114.444902174};
############ END DEBUG ############*/
test_input[39536:39543] = '{32'h41a6ebe6, 32'h42514b35, 32'h4249bc78, 32'hc28e8f25, 32'h41174d3b, 32'hc2c719fe, 32'h42b34bc4, 32'h42ae0838};
test_label[4942] = '{32'hc2c719fe};
test_output[4942] = '{32'h433d44aa};
/*############ DEBUG ############
test_input[39536:39543] = '{20.8651854441, 52.323445711, 50.4340520992, -71.2795781388, 9.45635525778, -99.5507629506, 89.647978969, 87.016050238};
test_label[4942] = '{-99.5507629506};
test_output[4942] = '{189.268211615};
############ END DEBUG ############*/
test_input[39544:39551] = '{32'hc15adee5, 32'hc10707e8, 32'h419f34ce, 32'hc1f75982, 32'hc11994fb, 32'hc12f41e9, 32'h429b8171, 32'h429b6b92};
test_label[4943] = '{32'h419f34ce};
test_output[4943] = '{32'h426a18a1};
/*############ DEBUG ############
test_input[39544:39551] = '{-13.6794173648, -8.43942979424, 19.9007839001, -30.9187055437, -9.59887262907, -10.9535917965, 77.7528159358, 77.7101020151};
test_label[4943] = '{19.9007839001};
test_output[4943] = '{58.5240502984};
############ END DEBUG ############*/
test_input[39552:39559] = '{32'hc25da5df, 32'h429692a9, 32'hc1c46b3a, 32'h42b42947, 32'hc023c234, 32'h428d08c0, 32'hc2b48ac1, 32'hc28a7e43};
test_label[4944] = '{32'h428d08c0};
test_output[4944] = '{32'h419c821e};
/*############ DEBUG ############
test_input[39552:39559] = '{-55.4119817708, 75.286446647, -24.552356069, 90.0806204078, -2.5587282637, 70.5170863098, -90.2710010735, -69.2466026702};
test_label[4944] = '{70.5170863098};
test_output[4944] = '{19.5635344769};
############ END DEBUG ############*/
test_input[39560:39567] = '{32'h425dd756, 32'h41dfea22, 32'h4286e87f, 32'hc28ce0e5, 32'hc263c45f, 32'hc081f149, 32'hc29927e7, 32'hc1eecd97};
test_label[4945] = '{32'hc263c45f};
test_output[4945] = '{32'h42f8cab0};
/*############ DEBUG ############
test_input[39560:39567] = '{55.4602896275, 27.9893233967, 67.4540966406, -70.439249236, -56.9417702205, -4.06070377728, -76.5779326983, -29.8503858719};
test_label[4945] = '{-56.9417702205};
test_output[4945] = '{124.395873043};
############ END DEBUG ############*/
test_input[39568:39575] = '{32'hc16ce071, 32'h42b06e7e, 32'hc2ad1eb9, 32'h3dcc096b, 32'h4222ee4b, 32'hc2068abc, 32'h42a4847b, 32'h42b31abf};
test_label[4946] = '{32'hc2ad1eb9};
test_output[4946] = '{32'h4330589a};
/*############ DEBUG ############
test_input[39568:39575] = '{-14.8047950354, 88.2158051935, -86.5600041272, 0.0996273378612, 40.7327070841, -33.6354822111, 82.2587508544, 89.552235536};
test_label[4946] = '{-86.5600041272};
test_output[4946] = '{176.34609523};
############ END DEBUG ############*/
test_input[39576:39583] = '{32'h4282af8b, 32'h424febe8, 32'h422017d6, 32'hc1e7e9cd, 32'hc2917035, 32'h419a50f1, 32'h41c584e6, 32'hc2c76703};
test_label[4947] = '{32'hc1e7e9cd};
test_output[4947] = '{32'h42bca9ff};
/*############ DEBUG ############
test_input[39576:39583] = '{65.3428588075, 51.9803764728, 40.023275944, -28.9891608563, -72.7191552794, 19.2895217529, 24.6898922039, -99.7011981787};
test_label[4947] = '{-28.9891608563};
test_output[4947] = '{94.3320212368};
############ END DEBUG ############*/
test_input[39584:39591] = '{32'hc2120248, 32'h42a688eb, 32'h425d8eba, 32'hc28bef28, 32'h42b69532, 32'hc27edd58, 32'h42a4f2c4, 32'hc011a485};
test_label[4948] = '{32'h42a4f2c4};
test_output[4948] = '{32'h410d1567};
/*############ DEBUG ############
test_input[39584:39591] = '{-36.5022283912, 83.2674175613, 55.3893813045, -69.967099736, 91.2913992984, -63.7161566758, 82.4741492178, -2.27566657963};
test_label[4948] = '{82.4741492178};
test_output[4948] = '{8.81772563607};
############ END DEBUG ############*/
test_input[39592:39599] = '{32'h4140b65d, 32'h421fa16d, 32'h412d465d, 32'hc1960274, 32'h4297471f, 32'hc053da73, 32'hc2737437, 32'hc2c660bc};
test_label[4949] = '{32'hc2737437};
test_output[4949] = '{32'h4308809d};
/*############ DEBUG ############
test_input[39592:39599] = '{12.0445226285, 39.9076422661, 10.8296783157, -18.7511978179, 75.6389089728, -3.31020815962, -60.8634911774, -99.1889365336};
test_label[4949] = '{-60.8634911774};
test_output[4949] = '{136.50240015};
############ END DEBUG ############*/
test_input[39600:39607] = '{32'h42ad3df6, 32'hc22b0002, 32'hc232496c, 32'h42831787, 32'h4206af6b, 32'h428e31af, 32'h4289c797, 32'hc29396b4};
test_label[4950] = '{32'h42831787};
test_output[4950] = '{32'h41a899bc};
/*############ DEBUG ############
test_input[39600:39607] = '{86.6210159334, -42.7500060435, -44.5717016589, 65.5459506764, 33.671307854, 71.0970346607, 68.8898243331, -73.7943436131};
test_label[4950] = '{65.5459506764};
test_output[4950] = '{21.0750654587};
############ END DEBUG ############*/
test_input[39608:39615] = '{32'hc1f06bf4, 32'h42897a90, 32'hc28a6714, 32'h40f5b617, 32'hc25086fb, 32'hc285ff65, 32'hbf8bfb48, 32'h42440959};
test_label[4951] = '{32'h40f5b617};
test_output[4951] = '{32'h42743e5d};
/*############ DEBUG ############
test_input[39608:39615] = '{-30.0527117785, 68.7393804347, -69.2013277354, 7.67847798815, -52.131818557, -66.9988144936, -1.09360604032, 49.0091280945};
test_label[4951] = '{7.67847798815};
test_output[4951] = '{61.0609024492};
############ END DEBUG ############*/
test_input[39616:39623] = '{32'hc2b14306, 32'hc1c887f2, 32'h41743e76, 32'h4229485a, 32'hc28e9d0a, 32'h42c3b10d, 32'hc055430c, 32'h42954bb6};
test_label[4952] = '{32'hc28e9d0a};
test_output[4952] = '{32'h4329270b};
/*############ DEBUG ############
test_input[39616:39623] = '{-88.6309080668, -25.0663803286, 15.2652489945, 42.3206575349, -71.3067148618, 97.8458043084, -3.33221716582, 74.6478711146};
test_label[4952] = '{-71.3067148618};
test_output[4952] = '{169.15251917};
############ END DEBUG ############*/
test_input[39624:39631] = '{32'hc229201a, 32'hc0b3d343, 32'hc2aafe98, 32'h426c1b46, 32'h425cba52, 32'hc2955b51, 32'h4221bfc9, 32'h4222f429};
test_label[4953] = '{32'hc2aafe98};
test_output[4953] = '{32'h43108b89};
/*############ DEBUG ############
test_input[39624:39631] = '{-42.2813476504, -5.61953870861, -85.4972571581, 59.0266342483, 55.1819543038, -74.6783488097, 40.4372919046, 40.7384386121};
test_label[4953] = '{-85.4972571581};
test_output[4953] = '{144.54505905};
############ END DEBUG ############*/
test_input[39632:39639] = '{32'h41974965, 32'h41a0db95, 32'hc119dea9, 32'h424717b2, 32'h42a6d59c, 32'hc211f347, 32'h401d283b, 32'h4142ae9f};
test_label[4954] = '{32'h41974965};
test_output[4954] = '{32'h42810343};
/*############ DEBUG ############
test_input[39632:39639] = '{18.9108368029, 20.1072178537, -9.61686085698, 49.7731387683, 83.4172081482, -36.487575496, 2.45558050665, 12.1676320214};
test_label[4954] = '{18.9108368029};
test_output[4954] = '{64.5063713454};
############ END DEBUG ############*/
test_input[39640:39647] = '{32'hc1596d07, 32'h42c7a2f9, 32'h42597d4d, 32'h42c22641, 32'hc2252438, 32'hc281d76d, 32'hc25f2438, 32'hc2b387e1};
test_label[4955] = '{32'h42c7a2f9};
test_output[4955] = '{32'h3d7f66d8};
/*############ DEBUG ############
test_input[39640:39647] = '{-13.5891183108, 99.8183064791, 54.372364858, 97.0747170113, -41.2853707235, -64.9207571697, -55.7853690483, -89.76538965};
test_label[4955] = '{99.8183064791};
test_output[4955] = '{0.0623539390322};
############ END DEBUG ############*/
test_input[39648:39655] = '{32'hc080c425, 32'hc2b3ad94, 32'h40e1f7a1, 32'hc2152aa9, 32'h41c6d501, 32'hc250d835, 32'hc1e8da9a, 32'h42c1a764};
test_label[4956] = '{32'hc2152aa9};
test_output[4956] = '{32'h43061e5c};
/*############ DEBUG ############
test_input[39648:39655] = '{-4.02394349047, -89.8390215573, 7.06147815212, -37.2916584503, 24.8540049344, -52.2111415332, -29.1067388544, 96.8269380463};
test_label[4956] = '{-37.2916584503};
test_output[4956] = '{134.118596497};
############ END DEBUG ############*/
test_input[39656:39663] = '{32'hc23149f6, 32'h421b8388, 32'h42a1505b, 32'hc2b6fd39, 32'hc2705234, 32'h405e1407, 32'hc2088115, 32'h425fe03a};
test_label[4957] = '{32'hc2088115};
test_output[4957] = '{32'h42e590e5};
/*############ DEBUG ############
test_input[39656:39663] = '{-44.3222269653, 38.878448126, 80.6569416868, -91.4945727389, -60.0802765423, 3.46997233126, -34.1260570774, 55.9689712962};
test_label[4957] = '{-34.1260570774};
test_output[4957] = '{114.782998764};
############ END DEBUG ############*/
test_input[39664:39671] = '{32'hc237a9c1, 32'h42229e7f, 32'h429496ae, 32'h41a80745, 32'h4201c488, 32'h3fb05eb2, 32'hc18477c4, 32'h42c6b79d};
test_label[4958] = '{32'h42229e7f};
test_output[4958] = '{32'h426ad0bc};
/*############ DEBUG ############
test_input[39664:39671] = '{-45.9157757198, 40.6547828372, 74.294297817, 21.0035491383, 32.4419244903, 1.3778899035, -16.5584799669, 99.3586232075};
test_label[4958] = '{40.6547828372};
test_output[4958] = '{58.7038403703};
############ END DEBUG ############*/
test_input[39672:39679] = '{32'h417dba0c, 32'hc2b65040, 32'hc2c1bd4d, 32'hc19b978b, 32'h3f5b4de9, 32'hc14ee87e, 32'h42a37d5b, 32'hc12ef52e};
test_label[4959] = '{32'hc19b978b};
test_output[4959] = '{32'h42ca633d};
/*############ DEBUG ############
test_input[39672:39679] = '{15.8579220304, -91.1567347294, -96.8697262576, -19.4489964419, 0.85665756844, -12.9317605167, 81.7448317052, -10.9348581689};
test_label[4959] = '{-19.4489964419};
test_output[4959] = '{101.193828147};
############ END DEBUG ############*/
test_input[39680:39687] = '{32'h426d64a3, 32'hc18b159c, 32'hc1120e73, 32'hc1becdca, 32'h41056da6, 32'hc20b7c97, 32'h41f45385, 32'h42027ed7};
test_label[4960] = '{32'h42027ed7};
test_output[4960] = '{32'h41d5cb97};
/*############ DEBUG ############
test_input[39680:39687] = '{59.3482780522, -17.3855519605, -9.1285281009, -23.8504827282, 8.33926979414, -34.8716686437, 30.5407805125, 32.6238681537};
test_label[4960] = '{32.6238681537};
test_output[4960] = '{26.7244098985};
############ END DEBUG ############*/
test_input[39688:39695] = '{32'hc13554fd, 32'hc2b444d8, 32'h42bcd652, 32'hc2789b66, 32'h429e1327, 32'h42bd62d2, 32'hc167941b, 32'hc22fc98d};
test_label[4961] = '{32'h42bcd652};
test_output[4961] = '{32'h3f56f91e};
/*############ DEBUG ############
test_input[39688:39695] = '{-11.3332486549, -90.1344596052, 94.4185961595, -62.15175659, 79.0374088759, 94.693011815, -14.4736583338, -43.9468287747};
test_label[4961] = '{94.4185961595};
test_output[4961] = '{0.839738705146};
############ END DEBUG ############*/
test_input[39696:39703] = '{32'hc1e9a1c1, 32'h421ba557, 32'h425cdcd2, 32'h42636f44, 32'hc2957e11, 32'h42047318, 32'h4200341b, 32'hc26de29b};
test_label[4962] = '{32'h425cdcd2};
test_output[4962] = '{32'h3fe8efbf};
/*############ DEBUG ############
test_input[39696:39703] = '{-29.2039819332, 38.9114638007, 55.215645189, 56.8586582605, -74.7462271006, 33.1123957832, 32.0508830736, -59.4712927566};
test_label[4962] = '{55.215645189};
test_output[4962] = '{1.8198164832};
############ END DEBUG ############*/
test_input[39704:39711] = '{32'hc269604f, 32'h420c7e2a, 32'hc1a1a9e9, 32'hc28d4e99, 32'h409f925b, 32'hc2551e57, 32'h3ef46077, 32'h423adb34};
test_label[4963] = '{32'h423adb34};
test_output[4963] = '{32'h371b317b};
/*############ DEBUG ############
test_input[39704:39711] = '{-58.3440513669, 35.123208484, -20.2079641756, -70.6535077558, 4.98661559059, -53.2796291158, 0.47729846286, 46.7140648336};
test_label[4963] = '{46.7140648336};
test_output[4963] = '{9.25024079602e-06};
############ END DEBUG ############*/
test_input[39712:39719] = '{32'h4298c4a7, 32'hbfbe01bd, 32'h419c35cd, 32'h42836c23, 32'hc2c533f1, 32'hc27c0bdf, 32'h42c45d8c, 32'hc2a4a5da};
test_label[4964] = '{32'hbfbe01bd};
test_output[4964] = '{32'h42c75593};
/*############ DEBUG ############
test_input[39712:39719] = '{76.3840895263, -1.48442800047, 19.526269481, 65.711207057, -98.6014459033, -63.0115926797, 98.1827053416, -82.3239308234};
test_label[4964] = '{-1.48442800047};
test_output[4964] = '{99.6671333424};
############ END DEBUG ############*/
test_input[39720:39727] = '{32'h419ff2d3, 32'hc2badb6f, 32'h425fe182, 32'h41edc248, 32'h41bc9567, 32'hc2325633, 32'h419d732d, 32'hc2928802};
test_label[4965] = '{32'h419ff2d3};
test_output[4965] = '{32'h420fe818};
/*############ DEBUG ############
test_input[39720:39727] = '{19.9935673502, -93.4285836524, 55.9702211859, 29.7198641436, 23.572950399, -44.5841782296, 19.6812374193, -73.2656409156};
test_label[4965] = '{19.9935673502};
test_output[4965] = '{35.9766538357};
############ END DEBUG ############*/
test_input[39728:39735] = '{32'h41f98717, 32'h429ec6c9, 32'hc1cd1b4c, 32'h41f1e35b, 32'hc24616b6, 32'hc27cd2ab, 32'h42487907, 32'hc22e5beb};
test_label[4966] = '{32'h429ec6c9};
test_output[4966] = '{32'h2a5a8000};
/*############ DEBUG ############
test_input[39728:39735] = '{31.1909614202, 79.388249648, -25.6383279953, 30.2360133712, -49.5221798821, -63.2057316901, 50.1181909538, -43.5897639657};
test_label[4966] = '{79.388249648};
test_output[4966] = '{1.94066984704e-13};
############ END DEBUG ############*/
test_input[39736:39743] = '{32'h429223db, 32'hc1f6781b, 32'h424f81f6, 32'h424c4df2, 32'hc2c7b08b, 32'hc25bc78d, 32'hc274f03c, 32'h429cbbe1};
test_label[4967] = '{32'h424f81f6};
test_output[4967] = '{32'h41d3f5d3};
/*############ DEBUG ############
test_input[39736:39743] = '{73.0700311254, -30.8086460681, 51.8769136763, 51.0761198468, -99.8448102098, -54.9448744943, -61.2346025717, 78.3669510464};
test_label[4967] = '{51.8769136763};
test_output[4967] = '{26.495031869};
############ END DEBUG ############*/
test_input[39744:39751] = '{32'h42c556d4, 32'h411c88a9, 32'hc2820f1b, 32'hc2135d74, 32'h429c0be1, 32'h42352855, 32'h4285e388, 32'h42235f89};
test_label[4968] = '{32'hc2820f1b};
test_output[4968] = '{32'h4323b2f7};
/*############ DEBUG ############
test_input[39744:39751] = '{98.6695827888, 9.783364459, -65.0295021358, -36.8412626983, 78.023204323, 45.2893883568, 66.9443995537, 40.8432945798};
test_label[4968] = '{-65.0295021358};
test_output[4968] = '{163.699084926};
############ END DEBUG ############*/
test_input[39752:39759] = '{32'h42b205b9, 32'hc1e86688, 32'hc2b9a90a, 32'hc2a47259, 32'h421d7116, 32'h424acf46, 32'h41963a16, 32'h428d8a72};
test_label[4969] = '{32'h42b205b9};
test_output[4969] = '{32'h324da8f4};
/*############ DEBUG ############
test_input[39752:39759] = '{89.0111804366, -29.0500646517, -92.8301519489, -82.2233339515, 39.3604366985, 50.7024168218, 18.7783615296, 70.7704005023};
test_label[4969] = '{89.0111804366};
test_output[4969] = '{1.19709861629e-08};
############ END DEBUG ############*/
test_input[39760:39767] = '{32'h41c30c35, 32'hc1fe7db9, 32'h42a23516, 32'h42673f8f, 32'hc1ed33fe, 32'h428a31a2, 32'hc242263b, 32'hc2c42f8a};
test_label[4970] = '{32'h42a23516};
test_output[4970] = '{32'h36ccc80a};
/*############ DEBUG ############
test_input[39760:39767] = '{24.3809605685, -31.8113875987, 81.1036852526, 57.8120680664, -29.6503865815, 69.0969393128, -48.537333613, -98.0928534667};
test_label[4970] = '{81.1036852526};
test_output[4970] = '{6.10296139629e-06};
############ END DEBUG ############*/
test_input[39768:39775] = '{32'h42ae02df, 32'hc1bfaad8, 32'hc1c5344a, 32'h425d6ca1, 32'hc20da433, 32'h424497f8, 32'h4113bbf6, 32'h425ee1b8};
test_label[4971] = '{32'h42ae02df};
test_output[4971] = '{32'h29458000};
/*############ DEBUG ############
test_input[39768:39775] = '{87.0056040994, -23.9584192097, -24.6505308495, 55.356083611, -35.410350347, 49.1484062303, 9.23338922968, 55.7204273038};
test_label[4971] = '{87.0056040994};
test_output[4971] = '{4.38538094727e-14};
############ END DEBUG ############*/
test_input[39776:39783] = '{32'hc198549c, 32'hc2683ddd, 32'hc249c5f2, 32'h4211343a, 32'hc218ac13, 32'h42089025, 32'h42662347, 32'hc251598a};
test_label[4972] = '{32'h4211343a};
test_output[4972] = '{32'h41a9de19};
/*############ DEBUG ############
test_input[39776:39783] = '{-19.0413129941, -58.06041473, -50.4433070593, 36.3010042851, -38.1680416874, 34.140767218, 57.5344503561, -52.3374394784};
test_label[4972] = '{36.3010042851};
test_output[4972] = '{21.2334460717};
############ END DEBUG ############*/
test_input[39784:39791] = '{32'h429f6007, 32'hc29fe626, 32'hc29b7f82, 32'hc2bd66ce, 32'hc09224e9, 32'h429194f8, 32'h42612854, 32'h42510113};
test_label[4973] = '{32'hc29fe626};
test_output[4973] = '{32'h431fa359};
/*############ DEBUG ############
test_input[39784:39791] = '{79.6875524649, -79.9495077502, -77.7490401826, -94.7007924177, -4.56700580015, 72.7909534371, 56.289381439, 52.2510480828};
test_label[4973] = '{-79.9495077502};
test_output[4973] = '{159.638070923};
############ END DEBUG ############*/
test_input[39792:39799] = '{32'h42204f03, 32'h42a0380d, 32'h423540cc, 32'hc1163ea8, 32'hc2b5465c, 32'hc285a179, 32'h426138c6, 32'h42565079};
test_label[4974] = '{32'h426138c6};
test_output[4974] = '{32'h41be6ea9};
/*############ DEBUG ############
test_input[39792:39799] = '{40.0771611701, 80.1094769029, 45.3132788299, -9.39029715253, -90.6374216703, -66.8153736644, 56.3054433298, 53.5785879425};
test_label[4974] = '{56.3054433298};
test_output[4974] = '{23.8040335732};
############ END DEBUG ############*/
test_input[39800:39807] = '{32'h4265a43c, 32'hc1e1344f, 32'hc2b7eebd, 32'h42a4b1b0, 32'hc2a85046, 32'hc287028d, 32'h42b13b62, 32'hc13747c6};
test_label[4975] = '{32'h4265a43c};
test_output[4975] = '{32'h41f9a8f0};
/*############ DEBUG ############
test_input[39800:39807] = '{57.410385315, -28.1505420848, -91.9662831774, 82.3470466652, -84.1567864338, -67.5049811818, 88.6159822913, -11.4550232268};
test_label[4975] = '{57.410385315};
test_output[4975] = '{31.2074894282};
############ END DEBUG ############*/
test_input[39808:39815] = '{32'hc18bb228, 32'hc1d5991f, 32'hc22302af, 32'hc1159225, 32'hc1ece0b8, 32'hc2bea7c3, 32'h42bf2ad3, 32'h42c40913};
test_label[4976] = '{32'h42c40913};
test_output[4976] = '{32'h3dac1ff8};
/*############ DEBUG ############
test_input[39808:39815] = '{-17.4619898784, -26.699766323, -40.7526215893, -9.34817939323, -29.609725824, -95.327660255, 95.5836425277, 98.0177242847};
test_label[4976] = '{98.0177242847};
test_output[4976] = '{0.0840453510214};
############ END DEBUG ############*/
test_input[39816:39823] = '{32'h41ec3856, 32'h425ed3f7, 32'h41a70711, 32'h42750eaf, 32'h424569f1, 32'h4236e400, 32'hc243bfba, 32'h42c4cbd7};
test_label[4977] = '{32'hc243bfba};
test_output[4977] = '{32'h431355da};
/*############ DEBUG ############
test_input[39816:39823] = '{29.5275080287, 55.7069987961, 20.8784502474, 61.264339842, 49.3534578583, 45.7226548408, -48.9372346365, 98.3981234207};
test_label[4977] = '{-48.9372346365};
test_output[4977] = '{147.335358057};
############ END DEBUG ############*/
test_input[39824:39831] = '{32'h425d157c, 32'hc0922c48, 32'hc20e6943, 32'h41068d33, 32'h42c3cd94, 32'hc2bd8bd3, 32'hc297142a, 32'hc252f6dc};
test_label[4978] = '{32'hc2bd8bd3};
test_output[4978] = '{32'h4340acb3};
/*############ DEBUG ############
test_input[39824:39831] = '{55.2709813112, -4.56790532129, -35.6027942122, 8.40947201705, 97.901519315, -94.7730919088, -75.5393793274, -52.7410734845};
test_label[4978] = '{-94.7730919088};
test_output[4978] = '{192.674611224};
############ END DEBUG ############*/
test_input[39832:39839] = '{32'hc2973f2a, 32'h427dc62e, 32'hc21da64d, 32'h41ef1d30, 32'hc2bd0e03, 32'hc2155b5c, 32'h4295d150, 32'h3fef8609};
test_label[4979] = '{32'h4295d150};
test_output[4979] = '{32'h372ff579};
/*############ DEBUG ############
test_input[39832:39839] = '{-75.6233708448, 63.443534689, -39.4124019702, 29.8892509617, -94.5273647992, -37.3392163688, 74.9088114799, 1.8712779403};
test_label[4979] = '{74.9088114799};
test_output[4979] = '{1.0487966193e-05};
############ END DEBUG ############*/
test_input[39840:39847] = '{32'hc2962ddc, 32'h42192127, 32'hc036a356, 32'h429ea551, 32'h415a345e, 32'h427ef8f2, 32'hc265a92f, 32'h4077954b};
test_label[4980] = '{32'h415a345e};
test_output[4980] = '{32'h42835ec5};
/*############ DEBUG ############
test_input[39840:39847] = '{-75.0895673546, 38.2823763005, -2.85371919532, 79.3228850715, 13.6377853799, 63.7431094011, -57.415218006, 3.8684871459};
test_label[4980] = '{13.6377853799};
test_output[4980] = '{65.685099863};
############ END DEBUG ############*/
test_input[39848:39855] = '{32'h42a07275, 32'h4256a266, 32'hc259807f, 32'h41cc3243, 32'h42a27918, 32'hc2b87a89, 32'hc16c4993, 32'hc28d4955};
test_label[4981] = '{32'h42a07275};
test_output[4981] = '{32'h3fa95002};
/*############ DEBUG ############
test_input[39848:39855] = '{80.2235472874, 53.6585935522, -54.3754839337, 25.5245415134, 81.2365093211, -92.2393271084, -14.767962855, -70.6432264973};
test_label[4981] = '{80.2235472874};
test_output[4981] = '{1.32275417728};
############ END DEBUG ############*/
test_input[39856:39863] = '{32'h4263f1a2, 32'hc248d772, 32'hc100f84e, 32'h422e267e, 32'hc1bd0517, 32'h42c7d005, 32'hc278d626, 32'hc0b88a19};
test_label[4982] = '{32'h42c7d005};
test_output[4982] = '{32'h80000000};
/*############ DEBUG ############
test_input[39856:39863] = '{56.9859696426, -50.2103954208, -8.06062146826, 43.5375904799, -23.6274853701, 99.9062860243, -62.2091286051, -5.76685739676};
test_label[4982] = '{99.9062860243};
test_output[4982] = '{-0.0};
############ END DEBUG ############*/
test_input[39864:39871] = '{32'hc29d2797, 32'hc28b839f, 32'h4021dc5e, 32'hc2bba623, 32'h41484243, 32'hc260aa94, 32'hc2656a2a, 32'h4090050b};
test_label[4983] = '{32'hc2656a2a};
test_output[4983] = '{32'h428bbd8f};
/*############ DEBUG ############
test_input[39864:39871] = '{-78.577321589, -69.7570719286, 2.52907512153, -93.8244820313, 12.5161768363, -56.1665786879, -57.3536772402, 4.50061553875};
test_label[4983] = '{-57.3536772402};
test_output[4983] = '{69.8702302778};
############ END DEBUG ############*/
test_input[39872:39879] = '{32'hc28142c5, 32'h428aed22, 32'hc2301828, 32'h42c1998e, 32'h423e300c, 32'h42bdd126, 32'h41b74e95, 32'hc280b483};
test_label[4984] = '{32'hc28142c5};
test_output[4984] = '{32'h43219222};
/*############ DEBUG ############
test_input[39872:39879] = '{-64.6304106492, 69.4631479122, -44.0235906793, 96.7999128069, 47.5469226125, 94.9084910746, 22.9133708837, -64.352563318};
test_label[4984] = '{-64.6304106492};
test_output[4984] = '{161.570830493};
############ END DEBUG ############*/
test_input[39880:39887] = '{32'hc27ef30a, 32'h4259c0dc, 32'hc2303c04, 32'h423394d3, 32'h41e2594a, 32'hc1814c11, 32'h421ae334, 32'hc2a42ed0};
test_label[4985] = '{32'hc2303c04};
test_output[4985] = '{32'h42c4fe79};
/*############ DEBUG ############
test_input[39880:39887] = '{-63.7373435727, 54.43834088, -44.0586074275, 44.8953359547, 28.2935984878, -16.162141062, 38.7218761859, -82.091432021};
test_label[4985] = '{-44.0586074275};
test_output[4985] = '{98.4970201554};
############ END DEBUG ############*/
test_input[39888:39895] = '{32'hc1f3de8f, 32'h4010a1c2, 32'h40130e37, 32'hc2b87c5e, 32'hc197ecd5, 32'hc049103c, 32'h400174c1, 32'hc1e0dfd1};
test_label[4986] = '{32'h4010a1c2};
test_output[4986] = '{32'h3f853ef3};
/*############ DEBUG ############
test_input[39888:39895] = '{-30.4836713938, 2.25987293789, 2.29774266291, -92.2429029742, -18.9906400955, -3.14161584275, 2.02275108316, -28.1092860972};
test_label[4986] = '{2.25987293789};
test_output[4986] = '{1.04098350595};
############ END DEBUG ############*/
test_input[39896:39903] = '{32'hc2405a25, 32'h42229715, 32'h3f89cfe2, 32'h4187610b, 32'h423c429b, 32'hc2b785f7, 32'hc285d8de, 32'hc23af4af};
test_label[4987] = '{32'h42229715};
test_output[4987] = '{32'h40cd698b};
/*############ DEBUG ############
test_input[39896:39903] = '{-48.0880310705, 40.6475418798, 1.07665659267, 16.9223836082, 47.0650441054, -91.7616517803, -66.9235684917, -46.7389476085};
test_label[4987] = '{40.6475418798};
test_output[4987] = '{6.41913362354};
############ END DEBUG ############*/
test_input[39904:39911] = '{32'hc2544d22, 32'h428eecb5, 32'h42946294, 32'hc0c1132e, 32'h429ef88e, 32'hc215e46d, 32'hc26c4b56, 32'hc2a01eb2};
test_label[4988] = '{32'h42946294};
test_output[4988] = '{32'h40a98b68};
/*############ DEBUG ############
test_input[39904:39911] = '{-53.0753261371, 71.4623219419, 74.1925349296, -6.0335914841, 79.4854618352, -37.4730715429, -59.0735702992, -80.0599537782};
test_label[4988] = '{74.1925349296};
test_output[4988] = '{5.29826743377};
############ END DEBUG ############*/
test_input[39912:39919] = '{32'hc179a471, 32'h41fd58cd, 32'h42b0bbe9, 32'h429c5b32, 32'hc2891848, 32'h4251c543, 32'h428a404e, 32'hc2204115};
test_label[4989] = '{32'h429c5b32};
test_output[4989] = '{32'h412305de};
/*############ DEBUG ############
test_input[39912:39919] = '{-15.6026471038, 31.6683588823, 88.3670086565, 78.1781134819, -68.5474277026, 52.4426374504, 69.1255926492, -40.0635575044};
test_label[4989] = '{78.1781134819};
test_output[4989] = '{10.1889327636};
############ END DEBUG ############*/
test_input[39920:39927] = '{32'h429b53ca, 32'h42b4f2fe, 32'h42a691b7, 32'hc295b99a, 32'hc2549e66, 32'hc21d061d, 32'h424914f7, 32'hc2addb8b};
test_label[4990] = '{32'hc2549e66};
test_output[4990] = '{32'h430fa14a};
/*############ DEBUG ############
test_input[39920:39927] = '{77.6636539624, 90.4745957919, 83.2845974268, -74.8625009886, -53.154684707, -39.2559703761, 50.2704746311, -86.9287924418};
test_label[4990] = '{-53.154684707};
test_output[4990] = '{143.630037034};
############ END DEBUG ############*/
test_input[39928:39935] = '{32'h42818426, 32'h429e9966, 32'hc23ca84a, 32'hc2c36abc, 32'hc2ab3116, 32'h4257beea, 32'h400a7135, 32'h420f054e};
test_label[4991] = '{32'hc2c36abc};
test_output[4991] = '{32'h43310211};
/*############ DEBUG ############
test_input[39928:39935] = '{64.7581041624, 79.2996085975, -47.1643430705, -97.7084661482, -85.5958729181, 53.936440453, 2.16315960591, 35.7551791946};
test_label[4991] = '{-97.7084661482};
test_output[4991] = '{177.00807523};
############ END DEBUG ############*/
test_input[39936:39943] = '{32'hc215df40, 32'h4280c690, 32'h42b8a140, 32'h42a8bf2e, 32'h41c9915e, 32'h4239cb03, 32'hc28f5832, 32'h426d56f9};
test_label[4992] = '{32'h41c9915e};
test_output[4992] = '{32'h42863d17};
/*############ DEBUG ############
test_input[39936:39943] = '{-37.4680187367, 64.3878159213, 92.3149385509, 84.3733992706, 25.1959796892, 46.4482549509, -71.6722547596, 59.3349352784};
test_label[4992] = '{25.1959796892};
test_output[4992] = '{67.1193144571};
############ END DEBUG ############*/
test_input[39944:39951] = '{32'hc1be62a7, 32'hc20a3112, 32'h413ab11d, 32'hc2b1c254, 32'h41fbc5e3, 32'h42285187, 32'h423be1a5, 32'h42024d81};
test_label[4993] = '{32'hc20a3112};
test_output[4993] = '{32'h42a30d31};
/*############ DEBUG ############
test_input[39944:39951] = '{-23.7981692384, -34.5479218467, 11.6682408622, -88.8795493831, 31.471623487, 42.0796172726, 46.9703573598, 32.5756863408};
test_label[4993] = '{-34.5479218467};
test_output[4993] = '{81.5257677018};
############ END DEBUG ############*/
test_input[39952:39959] = '{32'h404e1278, 32'h42ab3b53, 32'h422d2c37, 32'h428e4a76, 32'hc2c652a5, 32'hc2bea94f, 32'hc1ccaf9d, 32'hc280022a};
test_label[4994] = '{32'h404e1278};
test_output[4994] = '{32'h42a4cabf};
/*############ DEBUG ############
test_input[39952:39959] = '{3.2198771779, 85.6158656376, 43.2931774803, 71.1454325575, -99.1614161212, -95.3306806919, -25.5857487051, -64.0042288981};
test_label[4994] = '{3.2198771779};
test_output[4994] = '{82.3959889792};
############ END DEBUG ############*/
test_input[39960:39967] = '{32'h41c35a86, 32'h42625fe0, 32'hc1d87e7c, 32'hc245e3f1, 32'h42775040, 32'h42c785a9, 32'h41e66dbf, 32'h407923f9};
test_label[4995] = '{32'h42775040};
test_output[4995] = '{32'h4217bb11};
/*############ DEBUG ############
test_input[39960:39967] = '{24.4192016295, 56.593627724, -27.0617599564, -49.4725971649, 61.828371015, 99.7610547032, 28.8035875507, 3.89282050187};
test_label[4995] = '{61.828371015};
test_output[4995] = '{37.9326836882};
############ END DEBUG ############*/
test_input[39968:39975] = '{32'h42b1a71e, 32'hc072bda0, 32'h40d574c2, 32'h424d18b2, 32'hc288a694, 32'hc20fa952, 32'h40d5fbf3, 32'h410ad9a3};
test_label[4996] = '{32'hc072bda0};
test_output[4996] = '{32'h42b93d0b};
/*############ DEBUG ############
test_input[39968:39975] = '{88.8263973719, -3.7928237474, 6.67050264438, 51.2741178781, -68.3253442543, -35.9153508462, 6.68700529588, 8.67813380152};
test_label[4996] = '{-3.7928237474};
test_output[4996] = '{92.6192211193};
############ END DEBUG ############*/
test_input[39976:39983] = '{32'h413ee659, 32'hc2b9df63, 32'h40d52817, 32'hc2bd0c19, 32'h41c85308, 32'h425e1a6b, 32'hc2c2e497, 32'hc2c425a3};
test_label[4997] = '{32'hc2c425a3};
test_output[4997] = '{32'h4319996c};
/*############ DEBUG ############
test_input[39976:39983] = '{11.9312373853, -92.9363040173, 6.66114401703, -94.5236248658, 25.0405433346, 55.5257982142, -97.446465792, -98.0735066837};
test_label[4997] = '{-98.0735066837};
test_output[4997] = '{153.599304898};
############ END DEBUG ############*/
test_input[39984:39991] = '{32'h41f3176f, 32'hc29c858e, 32'h42393007, 32'h42bbc961, 32'hc2c6b98f, 32'h4268635a, 32'hc20c25c9, 32'hc21b4e7c};
test_label[4998] = '{32'h42bbc961};
test_output[4998] = '{32'h25c00000};
/*############ DEBUG ############
test_input[39984:39991] = '{30.3864430326, -78.2608503087, 46.2969035366, 93.8933157609, -99.3624228335, 58.0970214933, -35.0368983856, -38.8266435148};
test_label[4998] = '{93.8933157609};
test_output[4998] = '{3.33066907388e-16};
############ END DEBUG ############*/
test_input[39992:39999] = '{32'hc1dfa31a, 32'hc27743c0, 32'hc195b761, 32'hc1448b36, 32'h4240ba52, 32'hc1862780, 32'h424ce94c, 32'hc29e4ab9};
test_label[4999] = '{32'hc195b761};
test_output[4999] = '{32'h428bfa48};
/*############ DEBUG ############
test_input[39992:39999] = '{-27.9546402055, -61.8161612477, -18.714540975, -12.2839874825, 48.1819539869, -16.7692872784, 51.2278290214, -79.1459457869};
test_label[4999] = '{-18.714540975};
test_output[4999] = '{69.9888285701};
############ END DEBUG ############*/
end
`endif
