`ifndef SOFTMAX_WITH_LOSS_TEST_H
`define SOFTMAX_WITH_LOSS_TEST_H
reg [31:0] test_input [80];
reg [31:0] test_label [10];
reg [31:0] test_output [10];
initial begin
test_input[0:7] = '{32'h4288201d, 32'h41d39cf8, 32'hc1e4f432, 32'h41d6ec6b, 32'hc29c600d, 32'hc09a3152, 32'hc29cf9fe, 32'h419f3860};
test_label[0] = '{0};
test_output[0] = '{32'h80000000};
/*############ DEBUG ############
test_input[0:7] = '{68.0627243897, 26.4516441431, -28.6192357426, 26.8654379558, -78.1875956429, -4.81852042, -78.4882624073, 19.902526691};
test_label[0] = '{0};
test_output[0] = '{-0.0};
############ END DEBUG ############*/
test_input[8:15] = '{32'hc2402019, 32'hc26811eb, 32'h42b9e5cc, 32'h42beb82c, 32'hc22895a2, 32'hc2bdf9d2, 32'h429a97a2, 32'h429fa584};
test_label[1] = '{6};
test_output[1] = '{32'h41913228};
/*############ DEBUG ############
test_input[8:15] = '{-48.0313463489, -58.0174968351, 92.9488208643, 95.3597118986, -42.1461270734, -94.9879293892, 77.2961562969, 79.8232704965};
test_label[1] = '{6};
test_output[1] = '{18.1494906032};
############ END DEBUG ############*/
test_input[16:23] = '{32'hc233280d, 32'hc28c7a77, 32'hc18743cf, 32'hc2ae94f2, 32'hc216c300, 32'hc2b7df73, 32'hc2a9a3ac, 32'h41fd4754};
test_label[2] = '{3};
test_output[2] = '{32'h42ede6c7};
/*############ DEBUG ############
test_input[16:23] = '{-44.7891124572, -70.2391872381, -16.9081098649, -87.2909080821, -37.6904315227, -91.9364206336, -84.8196740048, 31.6598272412};
test_label[2] = '{3};
test_output[2] = '{118.950735323};
############ END DEBUG ############*/
test_input[24:31] = '{32'h4141befd, 32'hc23174df, 32'h42a2161d, 32'h42c6cd6e, 32'h42acb9c7, 32'hc24811e9, 32'hc2af5e99, 32'hc2ab183d};
test_label[3] = '{2};
test_output[3] = '{32'h4192dd46};
/*############ DEBUG ############
test_input[24:31] = '{12.1091278239, -44.3641310417, 81.0431914242, 99.4012327932, 86.3628454496, -50.0174920668, -87.684761512, -85.5473422729};
test_label[3] = '{2};
test_output[3] = '{18.3580435548};
############ END DEBUG ############*/
test_input[32:39] = '{32'hc0b7a985, 32'h42bf3ebc, 32'hc1e5e6ec, 32'h42537c46, 32'h40933d81, 32'hc26462cb, 32'h41e4b4a9, 32'hc27aea45};
test_label[4] = '{2};
test_output[4] = '{32'h42f8b877};
/*############ DEBUG ############
test_input[32:39] = '{-5.73944326795, 95.6225297759, -28.7377540815, 52.8713592167, 4.60125802615, -57.0964776424, 28.5882120589, -62.7287780161};
test_label[4] = '{2};
test_output[4] = '{124.360283857};
############ END DEBUG ############*/
test_input[40:47] = '{32'hc2744b4e, 32'h42a58376, 32'h4044f84c, 32'hc29c6845, 32'h41acea76, 32'h425edb71, 32'hc208c76b, 32'h421df151};
test_label[5] = '{6};
test_output[5] = '{32'h42e9e72c};
/*############ DEBUG ############
test_input[40:47] = '{-61.0735389726, 82.7567602399, 3.07765493955, -78.2036524884, 21.6144819406, 55.7142966748, -34.1947442746, 39.4856591549};
test_label[5] = '{6};
test_output[5] = '{116.951504514};
############ END DEBUG ############*/
test_input[48:55] = '{32'hc2682659, 32'hc2507dab, 32'h421d3d64, 32'hc2806c3d, 32'hc2303b8b, 32'h422c96e0, 32'hc00a9618, 32'hbfca27cd};
test_label[6] = '{4};
test_output[6] = '{32'h42ae7420};
/*############ DEBUG ############
test_input[48:55] = '{-58.037449063, -52.1227209817, 39.3099507374, -64.2114035012, -44.058147556, 43.1473404037, -2.16541110206, -1.57933963804};
test_label[6] = '{4};
test_output[6] = '{87.2268088262};
############ END DEBUG ############*/
test_input[56:63] = '{32'hc1718a4c, 32'h4157a2fb, 32'hc200178b, 32'hc29cacb2, 32'hc1fc45bb, 32'hc1c61848, 32'h41233c5a, 32'h423f7714};
test_label[7] = '{4};
test_output[7] = '{32'h429eccf9};
/*############ DEBUG ############
test_input[56:63] = '{-15.0962641339, 13.477290183, -32.0229895698, -78.3372927555, -31.5340474734, -24.7618567537, 10.2022342732, 47.8662873282};
test_label[7] = '{4};
test_output[7] = '{79.4003348016};
############ END DEBUG ############*/
test_input[64:71] = '{32'h42892dd3, 32'hc19b32e9, 32'hc161be9a, 32'h41df48b3, 32'hc1961ee6, 32'h4230804c, 32'h4167e7a1, 32'hc1e02870};
test_label[8] = '{6};
test_output[8] = '{32'h425861bd};
/*############ DEBUG ############
test_input[64:71] = '{68.5894982004, -19.3998580704, -14.1090331401, 27.9104970094, -18.7650876597, 44.1252898915, 14.4940503767, -28.019745733};
test_label[8] = '{6};
test_output[8] = '{54.0954478237};
############ END DEBUG ############*/
test_input[72:79] = '{32'h4271e905, 32'h42997c48, 32'hc294a410, 32'hc1da8428, 32'hc2b59848, 32'hc146127f, 32'hc23d7676, 32'h41c35e91};
test_label[9] = '{4};
test_output[9] = '{32'h43278a48};
/*############ DEBUG ############
test_input[72:79] = '{60.477556981, 76.7427362994, -74.3204378835, -27.3145300118, -90.7974266802, -12.3795155071, -47.3656831756, 24.4211745594};
test_label[9] = '{4};
test_output[9] = '{167.540163066};
############ END DEBUG ############*/
end
`endif
