../gen/afu_csr.vh